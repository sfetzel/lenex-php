<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="Breedy Badger" registration="LSV Tirol" version="11.42712">
    <CONTACT name="Breedy Badger" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" phone="+41 99 999 99 99" fax="+41 99 999 99 99" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Wien" name="Breedy Badger" name.en="3rd Int. Innsbrucker" course="LCM" deadline="2016-04-29" entrystartdate="2016-05-05" hostclub="" hostclub.url="" nation="AUT" organizer="" organizer.url="http://www.twv.at/" reservecount="2" result.url="http://www.schwimmverband-tirol.at/live/2016ibkmeet/index.html" startmethod="1" state="TI" timing="AUTOMATIC">
      <AGEDATE value="2016-05-07" type="YEAR" />
      <POOL name="Breedy Badger" lanemin="1" lanemax="8" />
      <POINTTABLE pointtableid="3005" name="Breedy Badger" version="2012" />
      <CONTACT city="Vienna" email="testfile@example.org" fax="+13 926315890234" name="Breedy Badger" phone="+43 (699) 10909741" street="Katzenbergerstrasse 2" zip="45879" />
      <QUALIFY from="2015-01-01" until="2016-04-29" />
      <SESSIONS>
        <SESSION date="2016-05-07" daytime="10:30" name="Breedy Badger" number="1" warmupfrom="09:30" warmupuntil="10:20">
          <EVENTS>
            <EVENT eventid="3649" daytime="13:47" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9785" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18195" />
                    <RANKING order="2" place="2" resultid="19060" />
                    <RANKING order="3" place="3" resultid="17294" />
                    <RANKING order="4" place="4" resultid="16616" />
                    <RANKING order="5" place="5" resultid="18433" />
                    <RANKING order="6" place="6" resultid="17288" />
                    <RANKING order="7" place="7" resultid="16640" />
                    <RANKING order="8" place="8" resultid="17300" />
                    <RANKING order="9" place="9" resultid="16599" />
                    <RANKING order="10" place="10" resultid="18255" />
                    <RANKING order="11" place="11" resultid="17282" />
                    <RANKING order="12" place="12" resultid="18442" />
                    <RANKING order="13" place="13" resultid="19225" />
                    <RANKING order="14" place="14" resultid="16938" />
                    <RANKING order="15" place="15" resultid="18714" />
                    <RANKING order="16" place="16" resultid="18204" />
                    <RANKING order="17" place="17" resultid="17499" />
                    <RANKING order="18" place="18" resultid="17874" />
                    <RANKING order="19" place="19" resultid="17908" />
                    <RANKING order="20" place="20" resultid="16933" />
                    <RANKING order="21" place="21" resultid="17414" />
                    <RANKING order="22" place="22" resultid="17949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9786" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16740" />
                    <RANKING order="2" place="2" resultid="17760" />
                    <RANKING order="3" place="3" resultid="18596" />
                    <RANKING order="4" place="4" resultid="17637" />
                    <RANKING order="5" place="5" resultid="16703" />
                    <RANKING order="6" place="6" resultid="19746" />
                    <RANKING order="7" place="7" resultid="17520" />
                    <RANKING order="8" place="8" resultid="17528" />
                    <RANKING order="9" place="9" resultid="17117" />
                    <RANKING order="10" place="10" resultid="17622" />
                    <RANKING order="11" place="11" resultid="18607" />
                    <RANKING order="12" place="12" resultid="18141" />
                    <RANKING order="13" place="13" resultid="17246" />
                    <RANKING order="14" place="14" resultid="17959" />
                    <RANKING order="15" place="15" resultid="16856" />
                    <RANKING order="16" place="16" resultid="17360" />
                    <RANKING order="17" place="17" resultid="17982" />
                    <RANKING order="18" place="18" resultid="16928" />
                    <RANKING order="19" place="19" resultid="18177" />
                    <RANKING order="20" place="20" resultid="16923" />
                    <RANKING order="21" place="21" resultid="19087" />
                    <RANKING order="22" place="22" resultid="16425" />
                    <RANKING order="23" place="23" resultid="19168" />
                    <RANKING order="24" place="-1" resultid="18773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9787" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18168" />
                    <RANKING order="2" place="2" resultid="18955" />
                    <RANKING order="3" place="3" resultid="18424" />
                    <RANKING order="4" place="4" resultid="17741" />
                    <RANKING order="5" place="5" resultid="17627" />
                    <RANKING order="6" place="6" resultid="18615" />
                    <RANKING order="7" place="7" resultid="16662" />
                    <RANKING order="8" place="8" resultid="17857" />
                    <RANKING order="9" place="9" resultid="18282" />
                    <RANKING order="10" place="10" resultid="17737" />
                    <RANKING order="11" place="11" resultid="17617" />
                    <RANKING order="12" place="12" resultid="17189" />
                    <RANKING order="13" place="13" resultid="17632" />
                    <RANKING order="14" place="14" resultid="17350" />
                    <RANKING order="15" place="15" resultid="18655" />
                    <RANKING order="16" place="16" resultid="16464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9788" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17468" />
                    <RANKING order="2" place="2" resultid="17687" />
                    <RANKING order="3" place="3" resultid="16731" />
                    <RANKING order="4" place="4" resultid="17097" />
                    <RANKING order="5" place="5" resultid="18647" />
                    <RANKING order="6" place="6" resultid="17697" />
                    <RANKING order="7" place="7" resultid="17226" />
                    <RANKING order="8" place="8" resultid="17394" />
                    <RANKING order="9" place="9" resultid="19109" />
                    <RANKING order="10" place="10" resultid="19719" />
                    <RANKING order="11" place="11" resultid="17334" />
                    <RANKING order="12" place="12" resultid="19114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9789" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9790" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19049" />
                    <RANKING order="2" place="2" resultid="18379" />
                    <RANKING order="3" place="3" resultid="19186" />
                    <RANKING order="4" place="4" resultid="17492" />
                    <RANKING order="5" place="5" resultid="19762" />
                    <RANKING order="6" place="6" resultid="19098" />
                    <RANKING order="7" place="7" resultid="18948" />
                    <RANKING order="8" place="8" resultid="16848" />
                    <RANKING order="9" place="9" resultid="19000" />
                    <RANKING order="10" place="10" resultid="17260" />
                    <RANKING order="11" place="11" resultid="19092" />
                    <RANKING order="12" place="12" resultid="17326" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19889" daytime="13:47" number="1" order="1" status="OFFICIAL" agegroupid="9790" />
                <HEAT heatid="19890" daytime="13:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19891" daytime="13:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19892" daytime="13:57" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19893" daytime="14:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19894" daytime="14:03" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19895" daytime="14:06" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19896" daytime="14:08" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19897" daytime="14:11" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19898" daytime="14:13" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19899" daytime="14:16" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3574" daytime="14:19" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3575" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18453" />
                    <RANKING order="2" place="2" resultid="19696" />
                    <RANKING order="3" place="3" resultid="16763" />
                    <RANKING order="4" place="4" resultid="19204" />
                    <RANKING order="5" place="5" resultid="19775" />
                    <RANKING order="6" place="6" resultid="18455" />
                    <RANKING order="7" place="7" resultid="19698" />
                    <RANKING order="8" place="8" resultid="19205" />
                    <RANKING order="9" place="9" resultid="18659" />
                    <RANKING order="10" place="10" resultid="18457" />
                    <RANKING order="11" place="11" resultid="19697" />
                    <RANKING order="12" place="12" resultid="17234" />
                    <RANKING order="13" place="13" resultid="19699" />
                    <RANKING order="14" place="14" resultid="16488" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20138" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20139" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3628" daytime="12:36" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9779" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17293" />
                    <RANKING order="2" place="2" resultid="19059" />
                    <RANKING order="3" place="3" resultid="17954" />
                    <RANKING order="4" place="4" resultid="18796" />
                    <RANKING order="5" place="5" resultid="16680" />
                    <RANKING order="6" place="6" resultid="19784" />
                    <RANKING order="7" place="7" resultid="17454" />
                    <RANKING order="8" place="8" resultid="18662" />
                    <RANKING order="9" place="9" resultid="16598" />
                    <RANKING order="10" place="10" resultid="18670" />
                    <RANKING order="11" place="11" resultid="18246" />
                    <RANKING order="12" place="12" resultid="17536" />
                    <RANKING order="13" place="13" resultid="19301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9780" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17429" />
                    <RANKING order="2" place="2" resultid="18618" />
                    <RANKING order="3" place="3" resultid="17602" />
                    <RANKING order="4" place="4" resultid="17755" />
                    <RANKING order="5" place="5" resultid="17750" />
                    <RANKING order="6" place="6" resultid="17532" />
                    <RANKING order="7" place="7" resultid="16671" />
                    <RANKING order="8" place="8" resultid="18911" />
                    <RANKING order="9" place="9" resultid="17368" />
                    <RANKING order="10" place="10" resultid="18186" />
                    <RANKING order="11" place="11" resultid="19126" />
                    <RANKING order="12" place="12" resultid="17902" />
                    <RANKING order="13" place="13" resultid="17153" />
                    <RANKING order="14" place="14" resultid="16781" />
                    <RANKING order="15" place="15" resultid="18000" />
                    <RANKING order="16" place="16" resultid="19167" />
                    <RANKING order="17" place="17" resultid="16710" />
                    <RANKING order="18" place="18" resultid="19272" />
                    <RANKING order="19" place="19" resultid="17672" />
                    <RANKING order="20" place="20" resultid="17667" />
                    <RANKING order="21" place="21" resultid="16424" />
                    <RANKING order="22" place="22" resultid="17587" />
                    <RANKING order="23" place="23" resultid="17386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9781" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17727" />
                    <RANKING order="2" place="2" resultid="17475" />
                    <RANKING order="3" place="3" resultid="18622" />
                    <RANKING order="4" place="4" resultid="17717" />
                    <RANKING order="5" place="5" resultid="17445" />
                    <RANKING order="6" place="6" resultid="18599" />
                    <RANKING order="7" place="7" resultid="16716" />
                    <RANKING order="8" place="8" resultid="19754" />
                    <RANKING order="9" place="9" resultid="19075" />
                    <RANKING order="10" place="10" resultid="16463" />
                    <RANKING order="11" place="10" resultid="18650" />
                    <RANKING order="12" place="12" resultid="17643" />
                    <RANKING order="13" place="13" resultid="17379" />
                    <RANKING order="14" place="14" resultid="18298" />
                    <RANKING order="15" place="15" resultid="18159" />
                    <RANKING order="16" place="16" resultid="18654" />
                    <RANKING order="17" place="-1" resultid="17722" />
                    <RANKING order="18" place="-1" resultid="18631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9782" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17692" />
                    <RANKING order="2" place="2" resultid="17702" />
                    <RANKING order="3" place="3" resultid="17437" />
                    <RANKING order="4" place="4" resultid="18646" />
                    <RANKING order="5" place="5" resultid="18983" />
                    <RANKING order="6" place="6" resultid="17022" />
                    <RANKING order="7" place="7" resultid="18132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9783" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17407" />
                    <RANKING order="2" place="2" resultid="17251" />
                    <RANKING order="3" place="3" resultid="17677" />
                    <RANKING order="4" place="4" resultid="19733" />
                    <RANKING order="5" place="5" resultid="17683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9784" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18611" />
                    <RANKING order="2" place="2" resultid="18938" />
                    <RANKING order="3" place="3" resultid="17325" />
                    <RANKING order="4" place="4" resultid="16420" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19864" daytime="12:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19865" daytime="12:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19866" daytime="12:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19867" daytime="12:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19868" daytime="12:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19869" daytime="12:46" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19870" daytime="12:47" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19871" daytime="12:49" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19872" daytime="12:51" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3621" daytime="12:14" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9763" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16864" />
                    <RANKING order="2" place="2" resultid="18890" />
                    <RANKING order="3" place="3" resultid="17896" />
                    <RANKING order="4" place="4" resultid="17162" />
                    <RANKING order="5" place="5" resultid="17842" />
                    <RANKING order="6" place="6" resultid="18776" />
                    <RANKING order="7" place="7" resultid="16589" />
                    <RANKING order="8" place="8" resultid="18820" />
                    <RANKING order="9" place="9" resultid="18698" />
                    <RANKING order="10" place="10" resultid="18231" />
                    <RANKING order="11" place="11" resultid="17198" />
                    <RANKING order="12" place="12" resultid="16580" />
                    <RANKING order="13" place="13" resultid="19042" />
                    <RANKING order="14" place="14" resultid="17504" />
                    <RANKING order="15" place="15" resultid="16958" />
                    <RANKING order="16" place="16" resultid="17524" />
                    <RANKING order="17" place="17" resultid="18690" />
                    <RANKING order="18" place="18" resultid="17884" />
                    <RANKING order="19" place="19" resultid="17662" />
                    <RANKING order="20" place="20" resultid="16967" />
                    <RANKING order="21" place="21" resultid="18018" />
                    <RANKING order="22" place="22" resultid="18678" />
                    <RANKING order="23" place="23" resultid="19003" />
                    <RANKING order="24" place="24" resultid="18964" />
                    <RANKING order="25" place="25" resultid="19289" />
                    <RANKING order="26" place="26" resultid="17861" />
                    <RANKING order="27" place="-1" resultid="18720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9764" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18850" />
                    <RANKING order="2" place="2" resultid="19055" />
                    <RANKING order="3" place="3" resultid="18290" />
                    <RANKING order="4" place="4" resultid="18551" />
                    <RANKING order="5" place="5" resultid="18566" />
                    <RANKING order="6" place="6" resultid="17799" />
                    <RANKING order="7" place="7" resultid="16790" />
                    <RANKING order="8" place="8" resultid="17126" />
                    <RANKING order="9" place="9" resultid="17171" />
                    <RANKING order="10" place="10" resultid="16648" />
                    <RANKING order="11" place="11" resultid="18554" />
                    <RANKING order="12" place="12" resultid="18033" />
                    <RANKING order="13" place="13" resultid="16432" />
                    <RANKING order="14" place="14" resultid="16687" />
                    <RANKING order="15" place="15" resultid="19027" />
                    <RANKING order="16" place="16" resultid="17375" />
                    <RANKING order="17" place="17" resultid="17820" />
                    <RANKING order="18" place="18" resultid="19120" />
                    <RANKING order="19" place="19" resultid="18509" />
                    <RANKING order="20" place="20" resultid="16822" />
                    <RANKING order="21" place="21" resultid="18498" />
                    <RANKING order="22" place="22" resultid="17048" />
                    <RANKING order="23" place="23" resultid="17013" />
                    <RANKING order="24" place="24" resultid="18213" />
                    <RANKING order="25" place="25" resultid="18495" />
                    <RANKING order="26" place="26" resultid="18014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9765" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17914" />
                    <RANKING order="2" place="2" resultid="18402" />
                    <RANKING order="3" place="3" resultid="18563" />
                    <RANKING order="4" place="4" resultid="18051" />
                    <RANKING order="5" place="5" resultid="17179" />
                    <RANKING order="6" place="6" resultid="17779" />
                    <RANKING order="7" place="7" resultid="18415" />
                    <RANKING order="8" place="8" resultid="18070" />
                    <RANKING order="9" place="9" resultid="18506" />
                    <RANKING order="10" place="10" resultid="18024" />
                    <RANKING order="11" place="11" resultid="17278" />
                    <RANKING order="12" place="12" resultid="17935" />
                    <RANKING order="13" place="13" resultid="18860" />
                    <RANKING order="14" place="14" resultid="18869" />
                    <RANKING order="15" place="15" resultid="17255" />
                    <RANKING order="16" place="16" resultid="16474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9766" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17144" />
                    <RANKING order="2" place="2" resultid="18578" />
                    <RANKING order="3" place="3" resultid="18900" />
                    <RANKING order="4" place="4" resultid="18037" />
                    <RANKING order="5" place="5" resultid="18106" />
                    <RANKING order="6" place="6" resultid="17273" />
                    <RANKING order="7" place="7" resultid="17044" />
                    <RANKING order="8" place="8" resultid="17003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9767" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18393" />
                    <RANKING order="2" place="2" resultid="18592" />
                    <RANKING order="3" place="3" resultid="18517" />
                    <RANKING order="4" place="4" resultid="16410" />
                    <RANKING order="5" place="5" resultid="18028" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19853" daytime="12:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19854" daytime="12:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19855" daytime="12:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19856" daytime="12:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19857" daytime="12:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19858" daytime="12:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19859" daytime="12:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19860" daytime="12:28" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19861" daytime="12:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19862" daytime="12:32" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19863" daytime="12:33" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3639" daytime="10:30" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3640" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17834" />
                    <RANKING order="2" place="2" resultid="19314" />
                    <RANKING order="3" place="3" resultid="16579" />
                    <RANKING order="4" place="4" resultid="18889" />
                    <RANKING order="5" place="5" resultid="17161" />
                    <RANKING order="6" place="6" resultid="16623" />
                    <RANKING order="7" place="7" resultid="16829" />
                    <RANKING order="8" place="8" resultid="17508" />
                    <RANKING order="9" place="9" resultid="17838" />
                    <RANKING order="10" place="10" resultid="19293" />
                    <RANKING order="11" place="11" resultid="16588" />
                    <RANKING order="12" place="12" resultid="18230" />
                    <RANKING order="13" place="13" resultid="18370" />
                    <RANKING order="14" place="14" resultid="17516" />
                    <RANKING order="15" place="15" resultid="17197" />
                    <RANKING order="16" place="16" resultid="17895" />
                    <RANKING order="17" place="17" resultid="17305" />
                    <RANKING order="18" place="18" resultid="17311" />
                    <RANKING order="19" place="19" resultid="16723" />
                    <RANKING order="20" place="20" resultid="18819" />
                    <RANKING order="21" place="21" resultid="17987" />
                    <RANKING order="22" place="22" resultid="18697" />
                    <RANKING order="23" place="23" resultid="16942" />
                    <RANKING order="24" place="24" resultid="18097" />
                    <RANKING order="25" place="25" resultid="18971" />
                    <RANKING order="26" place="26" resultid="19708" />
                    <RANKING order="27" place="27" resultid="18221" />
                    <RANKING order="28" place="28" resultid="18705" />
                    <RANKING order="29" place="29" resultid="19236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3642" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18570" />
                    <RANKING order="2" place="2" resultid="18849" />
                    <RANKING order="3" place="3" resultid="18337" />
                    <RANKING order="4" place="4" resultid="16607" />
                    <RANKING order="5" place="5" resultid="18550" />
                    <RANKING order="6" place="6" resultid="18346" />
                    <RANKING order="7" place="7" resultid="19054" />
                    <RANKING order="8" place="8" resultid="19007" />
                    <RANKING order="9" place="9" resultid="18289" />
                    <RANKING order="10" place="10" resultid="18088" />
                    <RANKING order="11" place="11" resultid="18988" />
                    <RANKING order="12" place="12" resultid="18150" />
                    <RANKING order="13" place="13" resultid="18529" />
                    <RANKING order="14" place="14" resultid="17264" />
                    <RANKING order="15" place="15" resultid="17105" />
                    <RANKING order="16" place="16" resultid="17125" />
                    <RANKING order="17" place="17" resultid="16647" />
                    <RANKING order="18" place="18" resultid="18542" />
                    <RANKING order="19" place="19" resultid="16789" />
                    <RANKING order="20" place="20" resultid="17825" />
                    <RANKING order="21" place="21" resultid="16753" />
                    <RANKING order="22" place="22" resultid="17170" />
                    <RANKING order="23" place="23" resultid="18032" />
                    <RANKING order="24" place="24" resultid="18355" />
                    <RANKING order="25" place="25" resultid="16686" />
                    <RANKING order="26" place="26" resultid="18272" />
                    <RANKING order="27" place="27" resultid="19014" />
                    <RANKING order="28" place="28" resultid="16451" />
                    <RANKING order="29" place="29" resultid="19026" />
                    <RANKING order="30" place="30" resultid="16430" />
                    <RANKING order="31" place="31" resultid="18013" />
                    <RANKING order="32" place="32" resultid="16813" />
                    <RANKING order="33" place="33" resultid="16821" />
                    <RANKING order="34" place="34" resultid="18212" />
                    <RANKING order="35" place="35" resultid="17993" />
                    <RANKING order="36" place="36" resultid="18385" />
                    <RANKING order="37" place="37" resultid="17373" />
                    <RANKING order="38" place="38" resultid="18043" />
                    <RANKING order="39" place="39" resultid="17920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3644" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18401" />
                    <RANKING order="2" place="2" resultid="17913" />
                    <RANKING order="3" place="3" resultid="16632" />
                    <RANKING order="4" place="4" resultid="18574" />
                    <RANKING order="5" place="5" resultid="18587" />
                    <RANKING order="6" place="6" resultid="18562" />
                    <RANKING order="7" place="7" resultid="18414" />
                    <RANKING order="8" place="8" resultid="17945" />
                    <RANKING order="9" place="9" resultid="18050" />
                    <RANKING order="10" place="10" resultid="18023" />
                    <RANKING order="11" place="11" resultid="17134" />
                    <RANKING order="12" place="12" resultid="17934" />
                    <RANKING order="13" place="13" resultid="16839" />
                    <RANKING order="14" place="14" resultid="18069" />
                    <RANKING order="15" place="15" resultid="19193" />
                    <RANKING order="16" place="16" resultid="18328" />
                    <RANKING order="17" place="17" resultid="17277" />
                    <RANKING order="18" place="18" resultid="17342" />
                    <RANKING order="19" place="18" resultid="18859" />
                    <RANKING order="20" place="20" resultid="16398" />
                    <RANKING order="21" place="21" resultid="16872" />
                    <RANKING order="22" place="22" resultid="17035" />
                    <RANKING order="23" place="23" resultid="18868" />
                    <RANKING order="24" place="24" resultid="16473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3645" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18524" />
                    <RANKING order="2" place="2" resultid="19727" />
                    <RANKING order="3" place="3" resultid="18239" />
                    <RANKING order="4" place="4" resultid="18319" />
                    <RANKING order="5" place="5" resultid="17143" />
                    <RANKING order="6" place="6" resultid="19722" />
                    <RANKING order="7" place="7" resultid="18105" />
                    <RANKING order="8" place="8" resultid="17774" />
                    <RANKING order="9" place="9" resultid="18899" />
                    <RANKING order="10" place="10" resultid="17053" />
                    <RANKING order="11" place="11" resultid="17272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3646" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18392" />
                    <RANKING order="2" place="2" resultid="18533" />
                    <RANKING order="3" place="3" resultid="17889" />
                    <RANKING order="4" place="4" resultid="18591" />
                    <RANKING order="5" place="5" resultid="19035" />
                    <RANKING order="6" place="6" resultid="16409" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19809" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19810" daytime="10:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19811" daytime="10:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19812" daytime="10:41" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19813" daytime="10:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19814" daytime="10:48" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19815" daytime="10:52" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19816" daytime="10:55" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19817" daytime="10:58" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19818" daytime="11:01" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19819" daytime="11:05" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19820" daytime="11:08" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19821" daytime="11:11" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19822" daytime="11:14" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3570" daytime="12:53" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9768" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16581" />
                    <RANKING order="2" place="2" resultid="16830" />
                    <RANKING order="3" place="3" resultid="16624" />
                    <RANKING order="4" place="4" resultid="17306" />
                    <RANKING order="5" place="5" resultid="18098" />
                    <RANKING order="6" place="6" resultid="19315" />
                    <RANKING order="7" place="7" resultid="16590" />
                    <RANKING order="8" place="8" resultid="18371" />
                    <RANKING order="9" place="9" resultid="17652" />
                    <RANKING order="10" place="10" resultid="19043" />
                    <RANKING order="11" place="11" resultid="19294" />
                    <RANKING order="12" place="12" resultid="16724" />
                    <RANKING order="13" place="13" resultid="17647" />
                    <RANKING order="14" place="14" resultid="18821" />
                    <RANKING order="15" place="15" resultid="17657" />
                    <RANKING order="16" place="16" resultid="17312" />
                    <RANKING order="17" place="17" resultid="18222" />
                    <RANKING order="18" place="18" resultid="17505" />
                    <RANKING order="19" place="19" resultid="19709" />
                    <RANKING order="20" place="20" resultid="18707" />
                    <RANKING order="21" place="21" resultid="16972" />
                    <RANKING order="22" place="22" resultid="18019" />
                    <RANKING order="23" place="23" resultid="16976" />
                    <RANKING order="24" place="24" resultid="18686" />
                    <RANKING order="25" place="25" resultid="16980" />
                    <RANKING order="26" place="26" resultid="19237" />
                    <RANKING order="27" place="27" resultid="18965" />
                    <RANKING order="28" place="28" resultid="19004" />
                    <RANKING order="29" place="29" resultid="16992" />
                    <RANKING order="30" place="30" resultid="16984" />
                    <RANKING order="31" place="31" resultid="16988" />
                    <RANKING order="32" place="32" resultid="18766" />
                    <RANKING order="33" place="-1" resultid="16996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9769" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18338" />
                    <RANKING order="2" place="2" resultid="16608" />
                    <RANKING order="3" place="3" resultid="17816" />
                    <RANKING order="4" place="4" resultid="19009" />
                    <RANKING order="5" place="5" resultid="18347" />
                    <RANKING order="6" place="6" resultid="17582" />
                    <RANKING order="7" place="7" resultid="18089" />
                    <RANKING order="8" place="8" resultid="18273" />
                    <RANKING order="9" place="9" resultid="17574" />
                    <RANKING order="10" place="10" resultid="18156" />
                    <RANKING order="11" place="11" resultid="18356" />
                    <RANKING order="12" place="12" resultid="17592" />
                    <RANKING order="13" place="13" resultid="18558" />
                    <RANKING order="14" place="14" resultid="17811" />
                    <RANKING order="15" place="15" resultid="16754" />
                    <RANKING order="16" place="16" resultid="18543" />
                    <RANKING order="17" place="17" resultid="17106" />
                    <RANKING order="18" place="18" resultid="18077" />
                    <RANKING order="19" place="19" resultid="18924" />
                    <RANKING order="20" place="20" resultid="17807" />
                    <RANKING order="21" place="21" resultid="18034" />
                    <RANKING order="22" place="22" resultid="16806" />
                    <RANKING order="23" place="23" resultid="16791" />
                    <RANKING order="24" place="24" resultid="19159" />
                    <RANKING order="25" place="25" resultid="17569" />
                    <RANKING order="26" place="26" resultid="16453" />
                    <RANKING order="27" place="27" resultid="16746" />
                    <RANKING order="28" place="28" resultid="19016" />
                    <RANKING order="29" place="29" resultid="18510" />
                    <RANKING order="30" place="30" resultid="18499" />
                    <RANKING order="31" place="31" resultid="18015" />
                    <RANKING order="32" place="32" resultid="16814" />
                    <RANKING order="33" place="33" resultid="17049" />
                    <RANKING order="34" place="34" resultid="18496" />
                    <RANKING order="35" place="35" resultid="17014" />
                    <RANKING order="36" place="36" resultid="18757" />
                    <RANKING order="37" place="-1" resultid="17976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9770" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16633" />
                    <RANKING order="2" place="2" resultid="17554" />
                    <RANKING order="3" place="3" resultid="17180" />
                    <RANKING order="4" place="4" resultid="19758" />
                    <RANKING order="5" place="5" resultid="17559" />
                    <RANKING order="6" place="6" resultid="18264" />
                    <RANKING order="7" place="7" resultid="16694" />
                    <RANKING order="8" place="8" resultid="18588" />
                    <RANKING order="9" place="9" resultid="18124" />
                    <RANKING order="10" place="10" resultid="17941" />
                    <RANKING order="11" place="11" resultid="18575" />
                    <RANKING order="12" place="12" resultid="17135" />
                    <RANKING order="13" place="13" resultid="19771" />
                    <RANKING order="14" place="14" resultid="17789" />
                    <RANKING order="15" place="15" resultid="18025" />
                    <RANKING order="16" place="16" resultid="16841" />
                    <RANKING order="17" place="17" resultid="17564" />
                    <RANKING order="18" place="18" resultid="18329" />
                    <RANKING order="19" place="19" resultid="18521" />
                    <RANKING order="20" place="20" resultid="17784" />
                    <RANKING order="21" place="21" resultid="17343" />
                    <RANKING order="22" place="22" resultid="18071" />
                    <RANKING order="23" place="23" resultid="17936" />
                    <RANKING order="24" place="24" resultid="18547" />
                    <RANKING order="25" place="25" resultid="16400" />
                    <RANKING order="26" place="26" resultid="17037" />
                    <RANKING order="27" place="27" resultid="17256" />
                    <RANKING order="28" place="28" resultid="16475" />
                    <RANKING order="29" place="29" resultid="18754" />
                    <RANKING order="30" place="30" resultid="18996" />
                    <RANKING order="31" place="31" resultid="18751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9771" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17846" />
                    <RANKING order="2" place="2" resultid="19729" />
                    <RANKING order="3" place="3" resultid="18320" />
                    <RANKING order="4" place="4" resultid="17549" />
                    <RANKING order="5" place="5" resultid="19723" />
                    <RANKING order="6" place="6" resultid="17851" />
                    <RANKING order="7" place="7" resultid="18579" />
                    <RANKING order="8" place="8" resultid="17055" />
                    <RANKING order="9" place="9" resultid="17004" />
                    <RANKING order="10" place="10" resultid="17009" />
                    <RANKING order="11" place="11" resultid="16442" />
                    <RANKING order="12" place="12" resultid="17045" />
                    <RANKING order="13" place="13" resultid="16404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9772" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18534" />
                    <RANKING order="2" place="2" resultid="17890" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19873" daytime="12:53" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19874" daytime="12:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19875" daytime="13:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19876" daytime="13:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19877" daytime="13:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19878" daytime="13:14" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19879" daytime="13:17" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19880" daytime="13:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19881" daytime="13:24" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19882" daytime="13:27" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19883" daytime="13:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19884" daytime="13:32" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19885" daytime="13:35" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19886" daytime="13:38" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="19887" daytime="13:41" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="19888" daytime="13:43" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="12820" daytime="14:32" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12821" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19692" />
                    <RANKING order="2" place="2" resultid="19201" />
                    <RANKING order="3" place="3" resultid="18450" />
                    <RANKING order="4" place="4" resultid="19200" />
                    <RANKING order="5" place="5" resultid="19693" />
                    <RANKING order="6" place="6" resultid="17465" />
                    <RANKING order="7" place="7" resultid="18660" />
                    <RANKING order="8" place="8" resultid="19694" />
                    <RANKING order="9" place="9" resultid="19774" />
                    <RANKING order="10" place="10" resultid="16761" />
                    <RANKING order="11" place="11" resultid="19695" />
                    <RANKING order="12" place="12" resultid="16487" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20140" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20141" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9711" daytime="11:17" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9713" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18194" />
                    <RANKING order="2" place="2" resultid="16615" />
                    <RANKING order="3" place="3" resultid="16639" />
                    <RANKING order="4" place="4" resultid="16679" />
                    <RANKING order="5" place="5" resultid="17287" />
                    <RANKING order="6" place="6" resultid="17953" />
                    <RANKING order="7" place="7" resultid="16597" />
                    <RANKING order="8" place="8" resultid="19224" />
                    <RANKING order="9" place="9" resultid="17299" />
                    <RANKING order="10" place="10" resultid="17281" />
                    <RANKING order="11" place="11" resultid="18669" />
                    <RANKING order="12" place="12" resultid="18432" />
                    <RANKING order="13" place="13" resultid="18245" />
                    <RANKING order="14" place="14" resultid="18310" />
                    <RANKING order="15" place="15" resultid="17948" />
                    <RANKING order="16" place="16" resultid="18203" />
                    <RANKING order="17" place="17" resultid="18441" />
                    <RANKING order="18" place="18" resultid="17413" />
                    <RANKING order="19" place="19" resultid="17453" />
                    <RANKING order="20" place="-1" resultid="19308" />
                    <RANKING order="21" place="-1" resultid="18661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9714" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16739" />
                    <RANKING order="2" place="2" resultid="17428" />
                    <RANKING order="3" place="3" resultid="17759" />
                    <RANKING order="4" place="4" resultid="16670" />
                    <RANKING order="5" place="5" resultid="17866" />
                    <RANKING order="6" place="6" resultid="16702" />
                    <RANKING order="7" place="7" resultid="17116" />
                    <RANKING order="8" place="8" resultid="17152" />
                    <RANKING order="9" place="9" resultid="18140" />
                    <RANKING order="10" place="10" resultid="16709" />
                    <RANKING order="11" place="11" resultid="17244" />
                    <RANKING order="12" place="12" resultid="17999" />
                    <RANKING order="13" place="13" resultid="17901" />
                    <RANKING order="14" place="14" resultid="17367" />
                    <RANKING order="15" place="15" resultid="19271" />
                    <RANKING order="16" place="16" resultid="17358" />
                    <RANKING order="17" place="17" resultid="18176" />
                    <RANKING order="18" place="18" resultid="17879" />
                    <RANKING order="19" place="19" resultid="16423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9715" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18167" />
                    <RANKING order="2" place="2" resultid="18626" />
                    <RANKING order="3" place="3" resultid="17712" />
                    <RANKING order="4" place="4" resultid="17206" />
                    <RANKING order="5" place="5" resultid="18423" />
                    <RANKING order="6" place="6" resultid="17856" />
                    <RANKING order="7" place="7" resultid="17612" />
                    <RANKING order="8" place="8" resultid="17607" />
                    <RANKING order="9" place="9" resultid="16715" />
                    <RANKING order="10" place="10" resultid="16661" />
                    <RANKING order="11" place="11" resultid="17597" />
                    <RANKING order="12" place="12" resultid="18634" />
                    <RANKING order="13" place="13" resultid="17349" />
                    <RANKING order="14" place="14" resultid="18281" />
                    <RANKING order="15" place="15" resultid="17642" />
                    <RANKING order="16" place="16" resultid="16462" />
                    <RANKING order="17" place="17" resultid="18158" />
                    <RANKING order="18" place="18" resultid="17378" />
                    <RANKING order="19" place="19" resultid="16483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9716" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18791" />
                    <RANKING order="2" place="2" resultid="17436" />
                    <RANKING order="3" place="3" resultid="17764" />
                    <RANKING order="4" place="4" resultid="16730" />
                    <RANKING order="5" place="5" resultid="19750" />
                    <RANKING order="6" place="6" resultid="18982" />
                    <RANKING order="7" place="7" resultid="17393" />
                    <RANKING order="8" place="8" resultid="17225" />
                    <RANKING order="9" place="9" resultid="17332" />
                    <RANKING order="10" place="10" resultid="19718" />
                    <RANKING order="11" place="11" resultid="17020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9717" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17406" />
                    <RANKING order="2" place="2" resultid="17250" />
                    <RANKING order="3" place="3" resultid="17682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9718" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19133" />
                    <RANKING order="2" place="2" resultid="19143" />
                    <RANKING order="3" place="3" resultid="18603" />
                    <RANKING order="4" place="4" resultid="18610" />
                    <RANKING order="5" place="5" resultid="18999" />
                    <RANKING order="6" place="6" resultid="17324" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19823" daytime="11:17" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19824" daytime="11:21" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19825" daytime="11:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19826" daytime="11:29" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19827" daytime="11:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19828" daytime="11:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19829" daytime="11:38" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19830" daytime="11:41" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19831" daytime="11:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19832" daytime="11:47" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3551" daytime="12:05" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9792" agemax="10" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18806" />
                    <RANKING order="2" place="2" resultid="19069" />
                    <RANKING order="3" place="3" resultid="19277" />
                    <RANKING order="4" place="4" resultid="17461" />
                    <RANKING order="5" place="5" resultid="17968" />
                    <RANKING order="6" place="6" resultid="17972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9773" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18713" />
                    <RANKING order="2" place="2" resultid="18254" />
                    <RANKING order="3" place="3" resultid="17873" />
                    <RANKING order="4" place="4" resultid="17540" />
                    <RANKING order="5" place="5" resultid="18311" />
                    <RANKING order="6" place="6" resultid="16937" />
                    <RANKING order="7" place="7" resultid="16932" />
                    <RANKING order="8" place="8" resultid="19788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9774" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17867" />
                    <RANKING order="2" place="2" resultid="19745" />
                    <RANKING order="3" place="3" resultid="18595" />
                    <RANKING order="4" place="4" resultid="17481" />
                    <RANKING order="5" place="5" resultid="18185" />
                    <RANKING order="6" place="6" resultid="16855" />
                    <RANKING order="7" place="7" resultid="17245" />
                    <RANKING order="8" place="8" resultid="16927" />
                    <RANKING order="9" place="9" resultid="16922" />
                    <RANKING order="10" place="10" resultid="17981" />
                    <RANKING order="11" place="11" resultid="19125" />
                    <RANKING order="12" place="12" resultid="19086" />
                    <RANKING order="13" place="13" resultid="17359" />
                    <RANKING order="14" place="14" resultid="19166" />
                    <RANKING order="15" place="15" resultid="17385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9775" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18954" />
                    <RANKING order="2" place="2" resultid="18614" />
                    <RANKING order="3" place="3" resultid="17474" />
                    <RANKING order="4" place="4" resultid="17707" />
                    <RANKING order="5" place="5" resultid="18627" />
                    <RANKING order="6" place="6" resultid="17207" />
                    <RANKING order="7" place="7" resultid="18635" />
                    <RANKING order="8" place="8" resultid="18630" />
                    <RANKING order="9" place="9" resultid="17188" />
                    <RANKING order="10" place="10" resultid="19074" />
                    <RANKING order="11" place="11" resultid="18297" />
                    <RANKING order="12" place="12" resultid="16484" />
                    <RANKING order="13" place="-1" resultid="17444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9776" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18363" />
                    <RANKING order="2" place="2" resultid="17421" />
                    <RANKING order="3" place="3" resultid="17096" />
                    <RANKING order="4" place="4" resultid="18642" />
                    <RANKING order="5" place="5" resultid="17333" />
                    <RANKING order="6" place="6" resultid="18131" />
                    <RANKING order="7" place="7" resultid="17021" />
                    <RANKING order="8" place="8" resultid="19108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9777" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9778" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17491" />
                    <RANKING order="2" place="2" resultid="19048" />
                    <RANKING order="3" place="3" resultid="16847" />
                    <RANKING order="4" place="4" resultid="19144" />
                    <RANKING order="5" place="5" resultid="19097" />
                    <RANKING order="6" place="6" resultid="17259" />
                    <RANKING order="7" place="7" resultid="18937" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19845" daytime="12:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19846" daytime="12:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19847" daytime="12:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19848" daytime="12:09" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19849" daytime="12:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19850" daytime="12:11" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19851" daytime="12:11" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19852" daytime="12:12" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3547" daytime="11:50" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9791" agemax="10" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18786" />
                    <RANKING order="2" place="2" resultid="17929" />
                    <RANKING order="3" place="3" resultid="19260" />
                    <RANKING order="4" place="4" resultid="18884" />
                    <RANKING order="5" place="5" resultid="18305" />
                    <RANKING order="6" place="6" resultid="19081" />
                    <RANKING order="7" place="7" resultid="19231" />
                    <RANKING order="8" place="8" resultid="17062" />
                    <RANKING order="9" place="9" resultid="19220" />
                    <RANKING order="10" place="10" resultid="17058" />
                    <RANKING order="11" place="11" resultid="18832" />
                    <RANKING order="12" place="12" resultid="17086" />
                    <RANKING order="13" place="13" resultid="19138" />
                    <RANKING order="14" place="14" resultid="18814" />
                    <RANKING order="15" place="15" resultid="19786" />
                    <RANKING order="16" place="16" resultid="17082" />
                    <RANKING order="17" place="17" resultid="19175" />
                    <RANKING order="18" place="18" resultid="17074" />
                    <RANKING order="19" place="19" resultid="17078" />
                    <RANKING order="20" place="20" resultid="18803" />
                    <RANKING order="21" place="21" resultid="17066" />
                    <RANKING order="22" place="22" resultid="17070" />
                    <RANKING order="23" place="23" resultid="18932" />
                    <RANKING order="24" place="24" resultid="18918" />
                    <RANKING order="25" place="25" resultid="17237" />
                    <RANKING order="26" place="26" resultid="18811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9758" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16863" />
                    <RANKING order="2" place="2" resultid="16943" />
                    <RANKING order="3" place="3" resultid="18685" />
                    <RANKING order="4" place="4" resultid="18677" />
                    <RANKING order="5" place="5" resultid="18706" />
                    <RANKING order="6" place="6" resultid="16957" />
                    <RANKING order="7" place="7" resultid="17512" />
                    <RANKING order="8" place="8" resultid="18689" />
                    <RANKING order="9" place="9" resultid="16979" />
                    <RANKING order="10" place="10" resultid="18021" />
                    <RANKING order="11" place="11" resultid="18963" />
                    <RANKING order="12" place="12" resultid="16995" />
                    <RANKING order="13" place="13" resultid="16975" />
                    <RANKING order="14" place="14" resultid="19002" />
                    <RANKING order="15" place="15" resultid="16983" />
                    <RANKING order="16" place="16" resultid="16971" />
                    <RANKING order="17" place="17" resultid="16991" />
                    <RANKING order="18" place="18" resultid="18765" />
                    <RANKING order="19" place="19" resultid="16987" />
                    <RANKING order="20" place="-1" resultid="18719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9759" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19151" />
                    <RANKING order="2" place="2" resultid="18923" />
                    <RANKING order="3" place="3" resultid="18076" />
                    <RANKING order="4" place="4" resultid="19158" />
                    <RANKING order="5" place="5" resultid="18513" />
                    <RANKING order="6" place="6" resultid="17265" />
                    <RANKING order="7" place="7" resultid="18530" />
                    <RANKING order="8" place="8" resultid="19015" />
                    <RANKING order="9" place="9" resultid="16805" />
                    <RANKING order="10" place="10" resultid="19008" />
                    <RANKING order="11" place="11" resultid="16452" />
                    <RANKING order="12" place="12" resultid="16431" />
                    <RANKING order="13" place="13" resultid="18386" />
                    <RANKING order="14" place="14" resultid="18583" />
                    <RANKING order="15" place="15" resultid="18044" />
                    <RANKING order="16" place="16" resultid="17374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9760" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17794" />
                    <RANKING order="2" place="2" resultid="16693" />
                    <RANKING order="3" place="3" resultid="19757" />
                    <RANKING order="4" place="4" resultid="18123" />
                    <RANKING order="5" place="5" resultid="18263" />
                    <RANKING order="6" place="6" resultid="18502" />
                    <RANKING order="7" place="7" resultid="19770" />
                    <RANKING order="8" place="8" resultid="18520" />
                    <RANKING order="9" place="9" resultid="16873" />
                    <RANKING order="10" place="10" resultid="19194" />
                    <RANKING order="11" place="11" resultid="16840" />
                    <RANKING order="12" place="12" resultid="18546" />
                    <RANKING order="13" place="13" resultid="16798" />
                    <RANKING order="14" place="14" resultid="17036" />
                    <RANKING order="15" place="15" resultid="16399" />
                    <RANKING order="16" place="16" resultid="18995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9761" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18525" />
                    <RANKING order="2" place="2" resultid="17544" />
                    <RANKING order="3" place="3" resultid="17769" />
                    <RANKING order="4" place="4" resultid="19737" />
                    <RANKING order="5" place="5" resultid="19728" />
                    <RANKING order="6" place="6" resultid="17008" />
                    <RANKING order="7" place="7" resultid="17054" />
                    <RANKING order="8" place="8" resultid="16441" />
                    <RANKING order="9" place="9" resultid="16403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9762" agemax="-1" agemin="19" name="Breedy Badger" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19833" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19834" daytime="11:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19835" daytime="11:53" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19836" daytime="11:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19837" daytime="11:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19838" daytime="11:57" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19839" daytime="11:58" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19840" daytime="11:59" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19841" daytime="12:00" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19842" daytime="12:01" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19843" daytime="12:02" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19844" daytime="12:03" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-05-07" daytime="14:45" name="Breedy Badger" number="2">
          <EVENTS>
            <EVENT eventid="15984" daytime="18:10" number="196" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15985" agemax="-1" agemin="-1" gender="F" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20157" />
                    <RANKING order="2" place="2" resultid="20188" />
                    <RANKING order="3" place="3" resultid="20171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15986" agemax="-1" agemin="-1" gender="M" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20228" />
                    <RANKING order="2" place="2" resultid="20231" />
                    <RANKING order="3" place="3" resultid="20214" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20130" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20131" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3505" daytime="16:36" gender="F" number="17" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9803" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16867" />
                    <RANKING order="2" place="2" resultid="16583" />
                    <RANKING order="3" place="3" resultid="16626" />
                    <RANKING order="4" place="4" resultid="18892" />
                    <RANKING order="5" place="5" resultid="18233" />
                    <RANKING order="6" place="6" resultid="16592" />
                    <RANKING order="7" place="7" resultid="17835" />
                    <RANKING order="8" place="8" resultid="17307" />
                    <RANKING order="9" place="9" resultid="17663" />
                    <RANKING order="10" place="10" resultid="18100" />
                    <RANKING order="11" place="11" resultid="17843" />
                    <RANKING order="12" place="12" resultid="19295" />
                    <RANKING order="13" place="13" resultid="17313" />
                    <RANKING order="14" place="14" resultid="18373" />
                    <RANKING order="15" place="15" resultid="16945" />
                    <RANKING order="16" place="16" resultid="18700" />
                    <RANKING order="17" place="17" resultid="18688" />
                    <RANKING order="18" place="18" resultid="18709" />
                    <RANKING order="19" place="19" resultid="19710" />
                    <RANKING order="20" place="20" resultid="18224" />
                    <RANKING order="21" place="21" resultid="18692" />
                    <RANKING order="22" place="22" resultid="18680" />
                    <RANKING order="23" place="23" resultid="17648" />
                    <RANKING order="24" place="24" resultid="17862" />
                    <RANKING order="25" place="-1" resultid="16725" />
                    <RANKING order="26" place="-1" resultid="18722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9804" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18853" />
                    <RANKING order="2" place="2" resultid="17583" />
                    <RANKING order="3" place="3" resultid="19153" />
                    <RANKING order="4" place="4" resultid="17266" />
                    <RANKING order="5" place="5" resultid="17812" />
                    <RANKING order="6" place="6" resultid="18340" />
                    <RANKING order="7" place="7" resultid="16610" />
                    <RANKING order="8" place="8" resultid="18079" />
                    <RANKING order="9" place="9" resultid="18531" />
                    <RANKING order="10" place="10" resultid="18926" />
                    <RANKING order="11" place="11" resultid="18091" />
                    <RANKING order="12" place="12" resultid="17826" />
                    <RANKING order="13" place="13" resultid="17571" />
                    <RANKING order="14" place="14" resultid="18358" />
                    <RANKING order="15" place="15" resultid="17808" />
                    <RANKING order="16" place="16" resultid="16756" />
                    <RANKING order="17" place="17" resultid="19161" />
                    <RANKING order="18" place="18" resultid="17108" />
                    <RANKING order="19" place="19" resultid="18515" />
                    <RANKING order="20" place="20" resultid="18275" />
                    <RANKING order="21" place="21" resultid="16748" />
                    <RANKING order="22" place="22" resultid="16808" />
                    <RANKING order="23" place="23" resultid="18215" />
                    <RANKING order="24" place="24" resultid="17994" />
                    <RANKING order="25" place="25" resultid="18585" />
                    <RANKING order="26" place="26" resultid="16435" />
                    <RANKING order="27" place="27" resultid="18046" />
                    <RANKING order="28" place="-1" resultid="19018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9805" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16696" />
                    <RANKING order="2" place="2" resultid="18266" />
                    <RANKING order="3" place="3" resultid="18126" />
                    <RANKING order="4" place="4" resultid="18589" />
                    <RANKING order="5" place="5" resultid="19760" />
                    <RANKING order="6" place="6" resultid="18504" />
                    <RANKING order="7" place="7" resultid="17790" />
                    <RANKING order="8" place="8" resultid="19773" />
                    <RANKING order="9" place="9" resultid="18522" />
                    <RANKING order="10" place="10" resultid="16875" />
                    <RANKING order="11" place="11" resultid="18331" />
                    <RANKING order="12" place="12" resultid="18862" />
                    <RANKING order="13" place="13" resultid="17345" />
                    <RANKING order="14" place="14" resultid="16800" />
                    <RANKING order="15" place="15" resultid="18870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9806" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18527" />
                    <RANKING order="2" place="2" resultid="17775" />
                    <RANKING order="3" place="3" resultid="19739" />
                    <RANKING order="4" place="4" resultid="17550" />
                    <RANKING order="5" place="5" resultid="18064" />
                    <RANKING order="6" place="6" resultid="17011" />
                    <RANKING order="7" place="7" resultid="16406" />
                    <RANKING order="8" place="-1" resultid="17852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9807" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19243" />
                    <RANKING order="2" place="2" resultid="16413" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19983" daytime="16:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19984" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19985" daytime="16:43" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19986" daytime="16:47" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19987" daytime="16:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19988" daytime="16:54" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19989" daytime="16:57" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19990" daytime="17:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19991" daytime="17:03" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19992" daytime="17:06" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19993" daytime="17:09" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="15921" daytime="17:55" number="191" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15971" agemax="-1" agemin="-1" gender="F" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20180" />
                    <RANKING order="2" place="2" resultid="20166" />
                    <RANKING order="3" place="3" resultid="20151" />
                    <RANKING order="4" place="4" resultid="20179" />
                    <RANKING order="5" place="5" resultid="20193" />
                    <RANKING order="6" place="6" resultid="20159" />
                    <RANKING order="7" place="7" resultid="20266" />
                    <RANKING order="8" place="8" resultid="20194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15928" agemax="-1" agemin="-1" gender="M" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20209" />
                    <RANKING order="2" place="2" resultid="20222" />
                    <RANKING order="3" place="3" resultid="20237" />
                    <RANKING order="4" place="4" resultid="20223" />
                    <RANKING order="5" place="5" resultid="20236" />
                    <RANKING order="6" place="6" resultid="20251" />
                    <RANKING order="7" place="7" resultid="20264" />
                    <RANKING order="8" place="8" resultid="20250" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20120" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20121" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="15987" daytime="18:13" number="197" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15988" agemax="-1" agemin="-1" gender="F" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20187" />
                    <RANKING order="2" place="2" resultid="20158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15989" agemax="-1" agemin="-1" gender="M" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20229" />
                    <RANKING order="2" place="2" resultid="20230" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20132" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20133" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="15972" daytime="17:58" number="192" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15973" agemax="-1" agemin="-1" gender="F" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20152" />
                    <RANKING order="2" place="2" resultid="20160" />
                    <RANKING order="3" place="3" resultid="20167" />
                    <RANKING order="4" place="4" resultid="20178" />
                    <RANKING order="5" place="5" resultid="20192" />
                    <RANKING order="6" place="6" resultid="20267" />
                    <RANKING order="7" place="7" resultid="20181" />
                    <RANKING order="8" place="-1" resultid="20203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15974" agemax="-1" agemin="-1" gender="M" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20224" />
                    <RANKING order="2" place="2" resultid="20210" />
                    <RANKING order="3" place="3" resultid="20238" />
                    <RANKING order="4" place="4" resultid="20221" />
                    <RANKING order="5" place="5" resultid="20252" />
                    <RANKING order="6" place="6" resultid="20235" />
                    <RANKING order="7" place="7" resultid="20263" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20122" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20123" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="15981" daytime="18:07" number="195" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15982" agemax="-1" agemin="-1" gender="F" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20189" />
                    <RANKING order="2" place="2" resultid="20156" />
                    <RANKING order="3" place="3" resultid="20170" />
                    <RANKING order="4" place="4" resultid="20163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15983" agemax="-1" agemin="-1" gender="M" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20232" />
                    <RANKING order="2" place="2" resultid="20213" />
                    <RANKING order="3" place="3" resultid="20227" />
                    <RANKING order="4" place="4" resultid="20241" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20128" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20129" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3538" daytime="14:45" gender="F" number="11" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9793" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16865" />
                    <RANKING order="2" place="2" resultid="18891" />
                    <RANKING order="3" place="3" resultid="17163" />
                    <RANKING order="4" place="4" resultid="17897" />
                    <RANKING order="5" place="5" resultid="16831" />
                    <RANKING order="6" place="6" resultid="18777" />
                    <RANKING order="7" place="7" resultid="18232" />
                    <RANKING order="8" place="8" resultid="17517" />
                    <RANKING order="9" place="9" resultid="18699" />
                    <RANKING order="10" place="10" resultid="17199" />
                    <RANKING order="11" place="11" resultid="18822" />
                    <RANKING order="12" place="12" resultid="18691" />
                    <RANKING order="13" place="13" resultid="17988" />
                    <RANKING order="14" place="14" resultid="16959" />
                    <RANKING order="15" place="15" resultid="16968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9794" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18851" />
                    <RANKING order="2" place="2" resultid="18291" />
                    <RANKING order="3" place="3" resultid="19056" />
                    <RANKING order="4" place="4" resultid="18552" />
                    <RANKING order="5" place="5" resultid="18567" />
                    <RANKING order="6" place="6" resultid="17127" />
                    <RANKING order="7" place="7" resultid="16792" />
                    <RANKING order="8" place="8" resultid="18555" />
                    <RANKING order="9" place="9" resultid="17172" />
                    <RANKING order="10" place="10" resultid="18149" />
                    <RANKING order="11" place="11" resultid="18090" />
                    <RANKING order="12" place="12" resultid="16649" />
                    <RANKING order="13" place="13" resultid="16688" />
                    <RANKING order="14" place="14" resultid="16433" />
                    <RANKING order="15" place="15" resultid="17821" />
                    <RANKING order="16" place="16" resultid="16815" />
                    <RANKING order="17" place="17" resultid="16823" />
                    <RANKING order="18" place="18" resultid="17050" />
                    <RANKING order="19" place="19" resultid="17015" />
                    <RANKING order="20" place="20" resultid="17977" />
                    <RANKING order="21" place="-1" resultid="19017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9795" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18403" />
                    <RANKING order="2" place="2" resultid="18564" />
                    <RANKING order="3" place="3" resultid="18416" />
                    <RANKING order="4" place="4" resultid="18052" />
                    <RANKING order="5" place="5" resultid="17181" />
                    <RANKING order="6" place="6" resultid="17279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9796" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17145" />
                    <RANKING order="2" place="2" resultid="18580" />
                    <RANKING order="3" place="3" resultid="17274" />
                    <RANKING order="4" place="4" resultid="17046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9797" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18394" />
                    <RANKING order="2" place="2" resultid="18593" />
                    <RANKING order="3" place="3" resultid="16411" />
                    <RANKING order="4" place="4" resultid="18029" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19904" daytime="14:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19905" daytime="14:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19906" daytime="14:53" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19907" daytime="14:57" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19908" daytime="15:01" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19909" daytime="15:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19910" daytime="15:08" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="15978" daytime="18:04" number="194" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15979" agemax="-1" agemin="-1" gender="F" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20155" />
                    <RANKING order="2" place="2" resultid="20169" />
                    <RANKING order="3" place="3" resultid="20190" />
                    <RANKING order="4" place="4" resultid="20162" />
                    <RANKING order="5" place="5" resultid="20176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15980" agemax="-1" agemin="-1" gender="M" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20233" />
                    <RANKING order="2" place="2" resultid="20212" />
                    <RANKING order="3" place="3" resultid="20226" />
                    <RANKING order="4" place="4" resultid="20240" />
                    <RANKING order="5" place="5" resultid="20254" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20126" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20127" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="20145" gender="F" number="190" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="20146" agemax="-1" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20149" />
                    <RANKING order="2" place="2" resultid="20150" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20148" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3562" daytime="16:23" gender="M" number="16" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9826" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19062" />
                    <RANKING order="2" place="2" resultid="16600" />
                    <RANKING order="3" place="3" resultid="18798" />
                    <RANKING order="4" place="4" resultid="18206" />
                    <RANKING order="5" place="5" resultid="18444" />
                    <RANKING order="6" place="6" resultid="16935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9827" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16741" />
                    <RANKING order="2" place="2" resultid="17756" />
                    <RANKING order="3" place="3" resultid="17623" />
                    <RANKING order="4" place="4" resultid="16673" />
                    <RANKING order="5" place="5" resultid="17521" />
                    <RANKING order="6" place="6" resultid="17745" />
                    <RANKING order="7" place="7" resultid="17668" />
                    <RANKING order="8" place="8" resultid="17673" />
                    <RANKING order="9" place="9" resultid="16930" />
                    <RANKING order="10" place="10" resultid="17880" />
                    <RANKING order="11" place="11" resultid="16428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9828" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17723" />
                    <RANKING order="2" place="2" resultid="18601" />
                    <RANKING order="3" place="3" resultid="17714" />
                    <RANKING order="4" place="4" resultid="17858" />
                    <RANKING order="5" place="5" resultid="18426" />
                    <RANKING order="6" place="6" resultid="17447" />
                    <RANKING order="7" place="7" resultid="16663" />
                    <RANKING order="8" place="8" resultid="18652" />
                    <RANKING order="9" place="9" resultid="17598" />
                    <RANKING order="10" place="10" resultid="18624" />
                    <RANKING order="11" place="11" resultid="17191" />
                    <RANKING order="12" place="12" resultid="17644" />
                    <RANKING order="13" place="13" resultid="16718" />
                    <RANKING order="14" place="14" resultid="18161" />
                    <RANKING order="15" place="15" resultid="16467" />
                    <RANKING order="16" place="16" resultid="16485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9829" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18365" />
                    <RANKING order="2" place="2" resultid="17765" />
                    <RANKING order="3" place="3" resultid="17099" />
                    <RANKING order="4" place="4" resultid="17698" />
                    <RANKING order="5" place="5" resultid="16732" />
                    <RANKING order="6" place="6" resultid="19752" />
                    <RANKING order="7" place="7" resultid="17439" />
                    <RANKING order="8" place="8" resultid="17396" />
                    <RANKING order="9" place="9" resultid="19720" />
                    <RANKING order="10" place="10" resultid="17336" />
                    <RANKING order="11" place="11" resultid="18134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9830" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9831" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18605" />
                    <RANKING order="2" place="2" resultid="17493" />
                    <RANKING order="3" place="3" resultid="18950" />
                    <RANKING order="4" place="4" resultid="19764" />
                    <RANKING order="5" place="5" resultid="19188" />
                    <RANKING order="6" place="6" resultid="19099" />
                    <RANKING order="7" place="7" resultid="16850" />
                    <RANKING order="8" place="8" resultid="18944" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19976" daytime="16:23" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19977" daytime="16:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19978" daytime="16:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19979" daytime="16:29" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19980" daytime="16:31" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19981" daytime="16:32" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19982" daytime="16:34" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="15975" daytime="18:01" number="193" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15976" agemax="-1" agemin="-1" gender="F" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20153" />
                    <RANKING order="2" place="2" resultid="20168" />
                    <RANKING order="3" place="3" resultid="20161" />
                    <RANKING order="4" place="4" resultid="20177" />
                    <RANKING order="5" place="5" resultid="20191" />
                    <RANKING order="6" place="6" resultid="20268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15977" agemax="-1" agemin="-1" gender="M" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20225" />
                    <RANKING order="2" place="2" resultid="20234" />
                    <RANKING order="3" place="3" resultid="20211" />
                    <RANKING order="4" place="4" resultid="20253" />
                    <RANKING order="5" place="5" resultid="20239" />
                    <RANKING order="6" place="6" resultid="20220" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20124" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20125" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3590" daytime="15:34" gender="F" number="13" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12822" agemax="10" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18787" />
                    <RANKING order="2" place="2" resultid="17930" />
                    <RANKING order="3" place="3" resultid="19261" />
                    <RANKING order="4" place="4" resultid="18885" />
                    <RANKING order="5" place="5" resultid="18306" />
                    <RANKING order="6" place="6" resultid="18833" />
                    <RANKING order="7" place="7" resultid="19082" />
                    <RANKING order="8" place="8" resultid="17060" />
                    <RANKING order="9" place="9" resultid="17076" />
                    <RANKING order="10" place="10" resultid="17064" />
                    <RANKING order="11" place="11" resultid="19232" />
                    <RANKING order="12" place="12" resultid="19176" />
                    <RANKING order="13" place="13" resultid="17084" />
                    <RANKING order="14" place="14" resultid="19221" />
                    <RANKING order="15" place="15" resultid="18459" />
                    <RANKING order="16" place="16" resultid="19139" />
                    <RANKING order="17" place="17" resultid="18783" />
                    <RANKING order="18" place="18" resultid="17072" />
                    <RANKING order="19" place="19" resultid="17087" />
                    <RANKING order="20" place="20" resultid="19787" />
                    <RANKING order="21" place="21" resultid="17238" />
                    <RANKING order="22" place="22" resultid="17068" />
                    <RANKING order="23" place="23" resultid="18815" />
                    <RANKING order="24" place="24" resultid="17080" />
                    <RANKING order="25" place="25" resultid="18804" />
                    <RANKING order="26" place="26" resultid="18933" />
                    <RANKING order="27" place="27" resultid="18919" />
                    <RANKING order="28" place="28" resultid="18812" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12823" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17509" />
                    <RANKING order="2" place="2" resultid="19316" />
                    <RANKING order="3" place="3" resultid="18099" />
                    <RANKING order="4" place="4" resultid="17200" />
                    <RANKING order="5" place="5" resultid="16944" />
                    <RANKING order="6" place="6" resultid="18778" />
                    <RANKING order="7" place="7" resultid="17513" />
                    <RANKING order="8" place="8" resultid="18708" />
                    <RANKING order="9" place="9" resultid="16960" />
                    <RANKING order="10" place="10" resultid="17525" />
                    <RANKING order="11" place="11" resultid="18223" />
                    <RANKING order="12" place="12" resultid="18020" />
                    <RANKING order="13" place="13" resultid="18059" />
                    <RANKING order="14" place="14" resultid="16969" />
                    <RANKING order="15" place="15" resultid="16981" />
                    <RANKING order="16" place="16" resultid="19005" />
                    <RANKING order="17" place="17" resultid="18966" />
                    <RANKING order="18" place="18" resultid="16977" />
                    <RANKING order="19" place="19" resultid="16973" />
                    <RANKING order="20" place="20" resultid="18679" />
                    <RANKING order="21" place="21" resultid="16997" />
                    <RANKING order="22" place="22" resultid="16985" />
                    <RANKING order="23" place="23" resultid="19238" />
                    <RANKING order="24" place="24" resultid="16993" />
                    <RANKING order="25" place="25" resultid="19290" />
                    <RANKING order="26" place="26" resultid="16989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12824" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18339" />
                    <RANKING order="2" place="2" resultid="18571" />
                    <RANKING order="3" place="3" resultid="16609" />
                    <RANKING order="4" place="4" resultid="18852" />
                    <RANKING order="5" place="5" resultid="18348" />
                    <RANKING order="6" place="6" resultid="18989" />
                    <RANKING order="7" place="7" resultid="18035" />
                    <RANKING order="8" place="8" resultid="18568" />
                    <RANKING order="9" place="9" resultid="16807" />
                    <RANKING order="10" place="10" resultid="18274" />
                    <RANKING order="11" place="11" resultid="18925" />
                    <RANKING order="12" place="12" resultid="19160" />
                    <RANKING order="13" place="13" resultid="18544" />
                    <RANKING order="14" place="14" resultid="19010" />
                    <RANKING order="15" place="15" resultid="18078" />
                    <RANKING order="16" place="16" resultid="18514" />
                    <RANKING order="17" place="17" resultid="17128" />
                    <RANKING order="18" place="18" resultid="18357" />
                    <RANKING order="19" place="19" resultid="18559" />
                    <RANKING order="20" place="20" resultid="16755" />
                    <RANKING order="21" place="21" resultid="17107" />
                    <RANKING order="22" place="22" resultid="17593" />
                    <RANKING order="23" place="23" resultid="16454" />
                    <RANKING order="24" place="24" resultid="18556" />
                    <RANKING order="25" place="25" resultid="18387" />
                    <RANKING order="26" place="26" resultid="17800" />
                    <RANKING order="27" place="27" resultid="16434" />
                    <RANKING order="28" place="28" resultid="17570" />
                    <RANKING order="29" place="28" resultid="19028" />
                    <RANKING order="30" place="30" resultid="18214" />
                    <RANKING order="31" place="31" resultid="16824" />
                    <RANKING order="32" place="32" resultid="16816" />
                    <RANKING order="33" place="33" resultid="18511" />
                    <RANKING order="34" place="34" resultid="18500" />
                    <RANKING order="35" place="35" resultid="17051" />
                    <RANKING order="36" place="36" resultid="18016" />
                    <RANKING order="37" place="37" resultid="17921" />
                    <RANKING order="38" place="38" resultid="17376" />
                    <RANKING order="39" place="39" resultid="18758" />
                    <RANKING order="40" place="40" resultid="18584" />
                    <RANKING order="41" place="41" resultid="18045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12825" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17915" />
                    <RANKING order="2" place="2" resultid="17560" />
                    <RANKING order="3" place="3" resultid="16634" />
                    <RANKING order="4" place="4" resultid="19759" />
                    <RANKING order="5" place="5" resultid="17795" />
                    <RANKING order="6" place="6" resultid="18404" />
                    <RANKING order="7" place="7" resultid="17942" />
                    <RANKING order="8" place="8" resultid="17182" />
                    <RANKING order="9" place="9" resultid="17780" />
                    <RANKING order="10" place="10" resultid="18026" />
                    <RANKING order="11" place="11" resultid="16695" />
                    <RANKING order="12" place="11" resultid="18503" />
                    <RANKING order="13" place="13" resultid="18265" />
                    <RANKING order="14" place="14" resultid="18125" />
                    <RANKING order="15" place="15" resultid="16842" />
                    <RANKING order="16" place="16" resultid="19772" />
                    <RANKING order="17" place="17" resultid="18072" />
                    <RANKING order="18" place="18" resultid="17344" />
                    <RANKING order="19" place="19" resultid="18330" />
                    <RANKING order="20" place="20" resultid="19195" />
                    <RANKING order="21" place="21" resultid="17257" />
                    <RANKING order="22" place="22" resultid="18548" />
                    <RANKING order="23" place="23" resultid="17280" />
                    <RANKING order="24" place="24" resultid="17937" />
                    <RANKING order="25" place="25" resultid="17785" />
                    <RANKING order="26" place="26" resultid="16874" />
                    <RANKING order="27" place="27" resultid="16401" />
                    <RANKING order="28" place="28" resultid="17038" />
                    <RANKING order="29" place="29" resultid="16476" />
                    <RANKING order="30" place="30" resultid="18755" />
                    <RANKING order="31" place="31" resultid="18997" />
                    <RANKING order="32" place="32" resultid="18752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12826" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18657" />
                    <RANKING order="2" place="2" resultid="17847" />
                    <RANKING order="3" place="3" resultid="19179" />
                    <RANKING order="4" place="4" resultid="19730" />
                    <RANKING order="5" place="5" resultid="19724" />
                    <RANKING order="6" place="6" resultid="18240" />
                    <RANKING order="7" place="7" resultid="18321" />
                    <RANKING order="8" place="8" resultid="17545" />
                    <RANKING order="9" place="9" resultid="18038" />
                    <RANKING order="10" place="10" resultid="19738" />
                    <RANKING order="11" place="11" resultid="18898" />
                    <RANKING order="12" place="12" resultid="18107" />
                    <RANKING order="13" place="13" resultid="17056" />
                    <RANKING order="14" place="14" resultid="18581" />
                    <RANKING order="15" place="15" resultid="18063" />
                    <RANKING order="16" place="16" resultid="17005" />
                    <RANKING order="17" place="17" resultid="17275" />
                    <RANKING order="18" place="18" resultid="16443" />
                    <RANKING order="19" place="19" resultid="17010" />
                    <RANKING order="20" place="20" resultid="16405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12827" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18395" />
                    <RANKING order="2" place="2" resultid="19715" />
                    <RANKING order="3" place="3" resultid="19242" />
                    <RANKING order="4" place="4" resultid="17891" />
                    <RANKING order="5" place="5" resultid="19036" />
                    <RANKING order="6" place="6" resultid="16412" />
                    <RANKING order="7" place="7" resultid="19149" />
                    <RANKING order="8" place="8" resultid="18518" />
                    <RANKING order="9" place="9" resultid="18030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12835" agemax="-1" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18657" />
                    <RANKING order="2" place="2" resultid="17915" />
                    <RANKING order="3" place="3" resultid="18395" />
                    <RANKING order="4" place="4" resultid="17847" />
                    <RANKING order="5" place="5" resultid="17560" />
                    <RANKING order="6" place="6" resultid="19715" />
                    <RANKING order="7" place="7" resultid="19179" />
                    <RANKING order="8" place="8" resultid="19242" />
                    <RANKING order="9" place="9" resultid="16634" />
                    <RANKING order="10" place="9" resultid="19730" />
                    <RANKING order="11" place="11" resultid="19724" />
                    <RANKING order="12" place="12" resultid="18240" />
                    <RANKING order="13" place="13" resultid="17891" />
                    <RANKING order="14" place="14" resultid="18339" />
                    <RANKING order="15" place="15" resultid="18571" />
                    <RANKING order="16" place="16" resultid="16609" />
                    <RANKING order="17" place="17" resultid="19759" />
                    <RANKING order="18" place="18" resultid="17795" />
                    <RANKING order="19" place="19" resultid="18404" />
                    <RANKING order="20" place="20" resultid="17942" />
                    <RANKING order="21" place="21" resultid="17182" />
                    <RANKING order="22" place="22" resultid="18321" />
                    <RANKING order="23" place="23" resultid="18852" />
                    <RANKING order="24" place="24" resultid="18348" />
                    <RANKING order="25" place="25" resultid="17780" />
                    <RANKING order="26" place="26" resultid="18026" />
                    <RANKING order="27" place="27" resultid="17545" />
                    <RANKING order="28" place="28" resultid="16695" />
                    <RANKING order="29" place="28" resultid="18503" />
                    <RANKING order="30" place="30" resultid="18989" />
                    <RANKING order="31" place="31" resultid="19036" />
                    <RANKING order="32" place="32" resultid="18038" />
                    <RANKING order="33" place="33" resultid="19738" />
                    <RANKING order="34" place="34" resultid="18265" />
                    <RANKING order="35" place="34" resultid="18898" />
                    <RANKING order="36" place="36" resultid="18035" />
                    <RANKING order="37" place="37" resultid="18125" />
                    <RANKING order="38" place="38" resultid="16842" />
                    <RANKING order="39" place="39" resultid="18568" />
                    <RANKING order="40" place="40" resultid="19772" />
                    <RANKING order="41" place="41" resultid="18072" />
                    <RANKING order="42" place="42" resultid="16807" />
                    <RANKING order="43" place="43" resultid="18274" />
                    <RANKING order="44" place="44" resultid="18925" />
                    <RANKING order="45" place="45" resultid="17344" />
                    <RANKING order="46" place="46" resultid="19160" />
                    <RANKING order="47" place="47" resultid="18544" />
                    <RANKING order="48" place="48" resultid="18107" />
                    <RANKING order="49" place="49" resultid="19010" />
                    <RANKING order="50" place="50" resultid="18330" />
                    <RANKING order="51" place="51" resultid="16412" />
                    <RANKING order="52" place="52" resultid="17056" />
                    <RANKING order="53" place="53" resultid="18581" />
                    <RANKING order="54" place="54" resultid="18078" />
                    <RANKING order="55" place="55" resultid="19195" />
                    <RANKING order="56" place="56" resultid="19149" />
                    <RANKING order="57" place="57" resultid="17509" />
                    <RANKING order="58" place="58" resultid="18514" />
                    <RANKING order="59" place="59" resultid="17128" />
                    <RANKING order="60" place="60" resultid="18357" />
                    <RANKING order="61" place="61" resultid="18559" />
                    <RANKING order="62" place="62" resultid="16755" />
                    <RANKING order="63" place="62" resultid="18518" />
                    <RANKING order="64" place="64" resultid="17107" />
                    <RANKING order="65" place="65" resultid="17593" />
                    <RANKING order="66" place="66" resultid="16454" />
                    <RANKING order="67" place="67" resultid="17257" />
                    <RANKING order="68" place="68" resultid="18548" />
                    <RANKING order="69" place="69" resultid="17280" />
                    <RANKING order="70" place="70" resultid="17937" />
                    <RANKING order="71" place="71" resultid="18556" />
                    <RANKING order="72" place="72" resultid="18030" />
                    <RANKING order="73" place="73" resultid="18387" />
                    <RANKING order="74" place="74" resultid="19316" />
                    <RANKING order="75" place="75" resultid="17800" />
                    <RANKING order="76" place="76" resultid="16434" />
                    <RANKING order="77" place="76" resultid="17785" />
                    <RANKING order="78" place="78" resultid="17570" />
                    <RANKING order="79" place="78" resultid="19028" />
                    <RANKING order="80" place="80" resultid="18214" />
                    <RANKING order="81" place="81" resultid="18063" />
                    <RANKING order="82" place="82" resultid="16874" />
                    <RANKING order="83" place="83" resultid="18787" />
                    <RANKING order="84" place="84" resultid="18099" />
                    <RANKING order="85" place="85" resultid="17200" />
                    <RANKING order="86" place="86" resultid="17930" />
                    <RANKING order="87" place="87" resultid="16401" />
                    <RANKING order="88" place="88" resultid="16824" />
                    <RANKING order="89" place="89" resultid="16816" />
                    <RANKING order="90" place="90" resultid="16944" />
                    <RANKING order="91" place="91" resultid="17005" />
                    <RANKING order="92" place="92" resultid="18511" />
                    <RANKING order="93" place="93" resultid="17038" />
                    <RANKING order="94" place="94" resultid="18778" />
                    <RANKING order="95" place="95" resultid="17275" />
                    <RANKING order="96" place="96" resultid="18500" />
                    <RANKING order="97" place="97" resultid="17513" />
                    <RANKING order="98" place="98" resultid="16443" />
                    <RANKING order="99" place="99" resultid="17051" />
                    <RANKING order="100" place="100" resultid="18708" />
                    <RANKING order="101" place="101" resultid="18016" />
                    <RANKING order="102" place="102" resultid="17921" />
                    <RANKING order="103" place="103" resultid="17376" />
                    <RANKING order="104" place="104" resultid="18758" />
                    <RANKING order="105" place="105" resultid="17010" />
                    <RANKING order="106" place="106" resultid="16960" />
                    <RANKING order="107" place="107" resultid="16476" />
                    <RANKING order="108" place="108" resultid="17525" />
                    <RANKING order="109" place="109" resultid="18223" />
                    <RANKING order="110" place="110" resultid="18755" />
                    <RANKING order="111" place="111" resultid="18020" />
                    <RANKING order="112" place="112" resultid="19261" />
                    <RANKING order="113" place="113" resultid="18584" />
                    <RANKING order="114" place="114" resultid="18045" />
                    <RANKING order="115" place="115" resultid="18059" />
                    <RANKING order="116" place="116" resultid="18885" />
                    <RANKING order="117" place="117" resultid="16405" />
                    <RANKING order="118" place="118" resultid="18306" />
                    <RANKING order="119" place="119" resultid="18997" />
                    <RANKING order="120" place="120" resultid="18833" />
                    <RANKING order="121" place="121" resultid="19082" />
                    <RANKING order="122" place="122" resultid="16969" />
                    <RANKING order="123" place="123" resultid="16981" />
                    <RANKING order="124" place="124" resultid="19005" />
                    <RANKING order="125" place="125" resultid="18966" />
                    <RANKING order="126" place="126" resultid="16977" />
                    <RANKING order="127" place="127" resultid="16973" />
                    <RANKING order="128" place="128" resultid="17060" />
                    <RANKING order="129" place="129" resultid="18679" />
                    <RANKING order="130" place="130" resultid="17076" />
                    <RANKING order="131" place="131" resultid="18752" />
                    <RANKING order="132" place="132" resultid="17064" />
                    <RANKING order="133" place="133" resultid="16997" />
                    <RANKING order="134" place="134" resultid="19232" />
                    <RANKING order="135" place="135" resultid="19176" />
                    <RANKING order="136" place="136" resultid="17084" />
                    <RANKING order="137" place="137" resultid="19221" />
                    <RANKING order="138" place="138" resultid="18459" />
                    <RANKING order="139" place="139" resultid="16985" />
                    <RANKING order="140" place="140" resultid="19139" />
                    <RANKING order="141" place="141" resultid="18783" />
                    <RANKING order="142" place="142" resultid="19238" />
                    <RANKING order="143" place="143" resultid="17072" />
                    <RANKING order="144" place="144" resultid="17087" />
                    <RANKING order="145" place="145" resultid="19787" />
                    <RANKING order="146" place="146" resultid="17238" />
                    <RANKING order="147" place="147" resultid="16993" />
                    <RANKING order="148" place="148" resultid="17068" />
                    <RANKING order="149" place="149" resultid="19290" />
                    <RANKING order="150" place="150" resultid="18815" />
                    <RANKING order="151" place="151" resultid="17080" />
                    <RANKING order="152" place="152" resultid="16989" />
                    <RANKING order="153" place="153" resultid="18804" />
                    <RANKING order="154" place="154" resultid="18933" />
                    <RANKING order="155" place="155" resultid="18919" />
                    <RANKING order="156" place="156" resultid="18812" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19917" daytime="15:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19918" daytime="15:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19919" daytime="15:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19920" daytime="15:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19921" daytime="15:39" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19922" daytime="15:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19923" daytime="15:41" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19924" daytime="15:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19925" daytime="15:43" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19926" daytime="15:44" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19927" daytime="15:45" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19928" daytime="15:46" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19929" daytime="15:47" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19930" daytime="15:47" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="19931" daytime="15:48" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="19932" daytime="15:49" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="19933" daytime="15:50" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="19934" daytime="15:51" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="19935" daytime="15:52" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="19936" daytime="15:52" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="19937" daytime="15:53" number="21" order="21" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3594" daytime="15:55" gender="M" number="14" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12828" agemax="10" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19070" />
                    <RANKING order="2" place="2" resultid="18807" />
                    <RANKING order="3" place="3" resultid="19278" />
                    <RANKING order="4" place="4" resultid="17462" />
                    <RANKING order="5" place="5" resultid="17488" />
                    <RANKING order="6" place="6" resultid="19305" />
                    <RANKING order="7" place="7" resultid="17969" />
                    <RANKING order="8" place="8" resultid="17973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12829" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18672" />
                    <RANKING order="2" place="2" resultid="17537" />
                    <RANKING order="3" place="3" resultid="18247" />
                    <RANKING order="4" place="4" resultid="19309" />
                    <RANKING order="5" place="5" resultid="19226" />
                    <RANKING order="6" place="6" resultid="18443" />
                    <RANKING order="7" place="7" resultid="16939" />
                    <RANKING order="8" place="8" resultid="18434" />
                    <RANKING order="9" place="9" resultid="18205" />
                    <RANKING order="10" place="10" resultid="18312" />
                    <RANKING order="11" place="11" resultid="17456" />
                    <RANKING order="12" place="12" resultid="16934" />
                    <RANKING order="13" place="13" resultid="19302" />
                    <RANKING order="14" place="14" resultid="17415" />
                    <RANKING order="15" place="15" resultid="19789" />
                    <RANKING order="16" place="-1" resultid="16617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12830" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18597" />
                    <RANKING order="2" place="2" resultid="17868" />
                    <RANKING order="3" place="3" resultid="17638" />
                    <RANKING order="4" place="4" resultid="17533" />
                    <RANKING order="5" place="5" resultid="17118" />
                    <RANKING order="6" place="6" resultid="17431" />
                    <RANKING order="7" place="7" resultid="19747" />
                    <RANKING order="8" place="8" resultid="18188" />
                    <RANKING order="9" place="9" resultid="18774" />
                    <RANKING order="10" place="10" resultid="18143" />
                    <RANKING order="11" place="11" resultid="17247" />
                    <RANKING order="12" place="12" resultid="16929" />
                    <RANKING order="13" place="13" resultid="17482" />
                    <RANKING order="14" place="14" resultid="18608" />
                    <RANKING order="15" place="15" resultid="18620" />
                    <RANKING order="16" place="16" resultid="18913" />
                    <RANKING order="17" place="17" resultid="17960" />
                    <RANKING order="18" place="18" resultid="19128" />
                    <RANKING order="19" place="19" resultid="18178" />
                    <RANKING order="20" place="20" resultid="16857" />
                    <RANKING order="21" place="21" resultid="17361" />
                    <RANKING order="22" place="22" resultid="16924" />
                    <RANKING order="23" place="23" resultid="19169" />
                    <RANKING order="24" place="24" resultid="19088" />
                    <RANKING order="25" place="25" resultid="17387" />
                    <RANKING order="26" place="26" resultid="16427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12831" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18956" />
                    <RANKING order="2" place="2" resultid="18425" />
                    <RANKING order="3" place="3" resultid="17476" />
                    <RANKING order="4" place="4" resultid="18616" />
                    <RANKING order="5" place="5" resultid="17732" />
                    <RANKING order="6" place="6" resultid="17628" />
                    <RANKING order="7" place="7" resultid="17613" />
                    <RANKING order="8" place="8" resultid="17713" />
                    <RANKING order="9" place="9" resultid="18169" />
                    <RANKING order="10" place="10" resultid="17209" />
                    <RANKING order="11" place="11" resultid="18600" />
                    <RANKING order="12" place="12" resultid="17446" />
                    <RANKING order="13" place="13" resultid="17351" />
                    <RANKING order="14" place="14" resultid="18283" />
                    <RANKING order="15" place="15" resultid="19755" />
                    <RANKING order="16" place="16" resultid="17618" />
                    <RANKING order="17" place="17" resultid="19076" />
                    <RANKING order="18" place="18" resultid="17608" />
                    <RANKING order="19" place="19" resultid="18651" />
                    <RANKING order="20" place="20" resultid="17190" />
                    <RANKING order="21" place="21" resultid="16466" />
                    <RANKING order="22" place="22" resultid="17633" />
                    <RANKING order="23" place="23" resultid="18632" />
                    <RANKING order="24" place="24" resultid="18299" />
                    <RANKING order="25" place="25" resultid="18160" />
                    <RANKING order="26" place="26" resultid="17380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12832" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18364" />
                    <RANKING order="2" place="2" resultid="17470" />
                    <RANKING order="3" place="3" resultid="17422" />
                    <RANKING order="4" place="4" resultid="19751" />
                    <RANKING order="5" place="5" resultid="17098" />
                    <RANKING order="6" place="6" resultid="17335" />
                    <RANKING order="7" place="7" resultid="19110" />
                    <RANKING order="8" place="8" resultid="18658" />
                    <RANKING order="9" place="9" resultid="18643" />
                    <RANKING order="10" place="9" resultid="19115" />
                    <RANKING order="11" place="11" resultid="17395" />
                    <RANKING order="12" place="12" resultid="18133" />
                    <RANKING order="13" place="13" resultid="17227" />
                    <RANKING order="14" place="14" resultid="17023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12833" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17408" />
                    <RANKING order="2" place="2" resultid="17678" />
                    <RANKING order="3" place="2" resultid="19768" />
                    <RANKING order="4" place="4" resultid="19735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12834" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19050" />
                    <RANKING order="2" place="2" resultid="19187" />
                    <RANKING order="3" place="3" resultid="19134" />
                    <RANKING order="4" place="4" resultid="18604" />
                    <RANKING order="5" place="5" resultid="19145" />
                    <RANKING order="6" place="6" resultid="18380" />
                    <RANKING order="7" place="7" resultid="18949" />
                    <RANKING order="8" place="8" resultid="19763" />
                    <RANKING order="9" place="9" resultid="16849" />
                    <RANKING order="10" place="10" resultid="18943" />
                    <RANKING order="11" place="11" resultid="19093" />
                    <RANKING order="12" place="12" resultid="17261" />
                    <RANKING order="13" place="13" resultid="18939" />
                    <RANKING order="14" place="14" resultid="17327" />
                    <RANKING order="15" place="15" resultid="19257" />
                    <RANKING order="16" place="16" resultid="16421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12852" agemax="-1" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19050" />
                    <RANKING order="2" place="2" resultid="19187" />
                    <RANKING order="3" place="3" resultid="19134" />
                    <RANKING order="4" place="4" resultid="18604" />
                    <RANKING order="5" place="5" resultid="19145" />
                    <RANKING order="6" place="6" resultid="18364" />
                    <RANKING order="7" place="7" resultid="18380" />
                    <RANKING order="8" place="8" resultid="18949" />
                    <RANKING order="9" place="9" resultid="18956" />
                    <RANKING order="10" place="10" resultid="17408" />
                    <RANKING order="11" place="11" resultid="19763" />
                    <RANKING order="12" place="12" resultid="16849" />
                    <RANKING order="13" place="13" resultid="18943" />
                    <RANKING order="14" place="14" resultid="17470" />
                    <RANKING order="15" place="15" resultid="18425" />
                    <RANKING order="16" place="16" resultid="17422" />
                    <RANKING order="17" place="17" resultid="19751" />
                    <RANKING order="18" place="18" resultid="17476" />
                    <RANKING order="19" place="19" resultid="18616" />
                    <RANKING order="20" place="20" resultid="17732" />
                    <RANKING order="21" place="21" resultid="17628" />
                    <RANKING order="22" place="22" resultid="17613" />
                    <RANKING order="23" place="23" resultid="17098" />
                    <RANKING order="24" place="24" resultid="17678" />
                    <RANKING order="25" place="24" resultid="17713" />
                    <RANKING order="26" place="24" resultid="19768" />
                    <RANKING order="27" place="27" resultid="18169" />
                    <RANKING order="28" place="28" resultid="19093" />
                    <RANKING order="29" place="29" resultid="17209" />
                    <RANKING order="30" place="30" resultid="18600" />
                    <RANKING order="31" place="31" resultid="17335" />
                    <RANKING order="32" place="31" resultid="17446" />
                    <RANKING order="33" place="33" resultid="17351" />
                    <RANKING order="34" place="34" resultid="18597" />
                    <RANKING order="35" place="35" resultid="19110" />
                    <RANKING order="36" place="36" resultid="18283" />
                    <RANKING order="37" place="37" resultid="18658" />
                    <RANKING order="38" place="38" resultid="18643" />
                    <RANKING order="39" place="38" resultid="19115" />
                    <RANKING order="40" place="40" resultid="17395" />
                    <RANKING order="41" place="41" resultid="17261" />
                    <RANKING order="42" place="42" resultid="17868" />
                    <RANKING order="43" place="43" resultid="18939" />
                    <RANKING order="44" place="43" resultid="19755" />
                    <RANKING order="45" place="45" resultid="18133" />
                    <RANKING order="46" place="46" resultid="17227" />
                    <RANKING order="47" place="47" resultid="17638" />
                    <RANKING order="48" place="48" resultid="17618" />
                    <RANKING order="49" place="49" resultid="17533" />
                    <RANKING order="50" place="50" resultid="17327" />
                    <RANKING order="51" place="51" resultid="19076" />
                    <RANKING order="52" place="52" resultid="17023" />
                    <RANKING order="53" place="53" resultid="19735" />
                    <RANKING order="54" place="54" resultid="17608" />
                    <RANKING order="55" place="55" resultid="18651" />
                    <RANKING order="56" place="56" resultid="17190" />
                    <RANKING order="57" place="57" resultid="16466" />
                    <RANKING order="58" place="58" resultid="17633" />
                    <RANKING order="59" place="59" resultid="17118" />
                    <RANKING order="60" place="60" resultid="17431" />
                    <RANKING order="61" place="61" resultid="18632" />
                    <RANKING order="62" place="62" resultid="19747" />
                    <RANKING order="63" place="63" resultid="18299" />
                    <RANKING order="64" place="64" resultid="18160" />
                    <RANKING order="65" place="65" resultid="18188" />
                    <RANKING order="66" place="66" resultid="17380" />
                    <RANKING order="67" place="67" resultid="18774" />
                    <RANKING order="68" place="68" resultid="18143" />
                    <RANKING order="69" place="69" resultid="17247" />
                    <RANKING order="70" place="70" resultid="16929" />
                    <RANKING order="71" place="71" resultid="17482" />
                    <RANKING order="72" place="72" resultid="18608" />
                    <RANKING order="73" place="73" resultid="18620" />
                    <RANKING order="74" place="74" resultid="18913" />
                    <RANKING order="75" place="75" resultid="17960" />
                    <RANKING order="76" place="76" resultid="19128" />
                    <RANKING order="77" place="77" resultid="19257" />
                    <RANKING order="78" place="78" resultid="18178" />
                    <RANKING order="79" place="79" resultid="18672" />
                    <RANKING order="80" place="80" resultid="16857" />
                    <RANKING order="81" place="81" resultid="17361" />
                    <RANKING order="82" place="82" resultid="16924" />
                    <RANKING order="83" place="83" resultid="17537" />
                    <RANKING order="84" place="84" resultid="18247" />
                    <RANKING order="85" place="85" resultid="16421" />
                    <RANKING order="86" place="86" resultid="19309" />
                    <RANKING order="87" place="87" resultid="19226" />
                    <RANKING order="88" place="88" resultid="18443" />
                    <RANKING order="89" place="88" resultid="19169" />
                    <RANKING order="90" place="90" resultid="16939" />
                    <RANKING order="91" place="91" resultid="18434" />
                    <RANKING order="92" place="92" resultid="19088" />
                    <RANKING order="93" place="93" resultid="18205" />
                    <RANKING order="94" place="94" resultid="18312" />
                    <RANKING order="95" place="95" resultid="17456" />
                    <RANKING order="96" place="96" resultid="19070" />
                    <RANKING order="97" place="97" resultid="18807" />
                    <RANKING order="98" place="98" resultid="16934" />
                    <RANKING order="99" place="99" resultid="19278" />
                    <RANKING order="100" place="100" resultid="17387" />
                    <RANKING order="101" place="101" resultid="16427" />
                    <RANKING order="102" place="102" resultid="19302" />
                    <RANKING order="103" place="103" resultid="17415" />
                    <RANKING order="104" place="104" resultid="17462" />
                    <RANKING order="105" place="105" resultid="17488" />
                    <RANKING order="106" place="106" resultid="19789" />
                    <RANKING order="107" place="107" resultid="19305" />
                    <RANKING order="108" place="108" resultid="17969" />
                    <RANKING order="109" place="109" resultid="17973" />
                    <RANKING order="110" place="-1" resultid="16617" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19945" daytime="15:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19946" daytime="15:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19947" daytime="15:57" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19948" daytime="15:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19949" daytime="15:59" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19950" daytime="16:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19951" daytime="16:01" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19952" daytime="16:02" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19953" daytime="16:03" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19954" daytime="16:04" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19955" daytime="16:04" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19956" daytime="16:05" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19957" daytime="16:06" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19958" daytime="16:07" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="19959" daytime="16:08" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3555" daytime="16:09" gender="F" number="15" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9798" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16866" />
                    <RANKING order="2" place="2" resultid="16582" />
                    <RANKING order="3" place="3" resultid="17830" />
                    <RANKING order="4" place="4" resultid="19317" />
                    <RANKING order="5" place="5" resultid="17653" />
                    <RANKING order="6" place="6" resultid="17164" />
                    <RANKING order="7" place="7" resultid="16591" />
                    <RANKING order="8" place="8" resultid="16625" />
                    <RANKING order="9" place="9" resultid="18372" />
                    <RANKING order="10" place="10" resultid="19044" />
                    <RANKING order="11" place="11" resultid="18972" />
                    <RANKING order="12" place="12" resultid="17658" />
                    <RANKING order="13" place="13" resultid="17989" />
                    <RANKING order="14" place="14" resultid="16832" />
                    <RANKING order="15" place="15" resultid="18687" />
                    <RANKING order="16" place="16" resultid="17885" />
                    <RANKING order="17" place="-1" resultid="18721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9799" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18572" />
                    <RANKING order="2" place="2" resultid="19152" />
                    <RANKING order="3" place="3" resultid="18990" />
                    <RANKING order="4" place="4" resultid="18560" />
                    <RANKING order="5" place="5" resultid="19057" />
                    <RANKING order="6" place="6" resultid="17575" />
                    <RANKING order="7" place="7" resultid="18151" />
                    <RANKING order="8" place="8" resultid="18349" />
                    <RANKING order="9" place="9" resultid="18292" />
                    <RANKING order="10" place="10" resultid="17173" />
                    <RANKING order="11" place="11" resultid="16747" />
                    <RANKING order="12" place="12" resultid="16793" />
                    <RANKING order="13" place="13" resultid="19029" />
                    <RANKING order="14" place="14" resultid="16455" />
                    <RANKING order="15" place="15" resultid="19121" />
                    <RANKING order="16" place="-1" resultid="17803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9800" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16635" />
                    <RANKING order="2" place="2" resultid="18576" />
                    <RANKING order="3" place="3" resultid="17555" />
                    <RANKING order="4" place="4" resultid="16843" />
                    <RANKING order="5" place="5" resultid="18053" />
                    <RANKING order="6" place="6" resultid="18507" />
                    <RANKING order="7" place="7" resultid="18417" />
                    <RANKING order="8" place="8" resultid="17565" />
                    <RANKING order="9" place="9" resultid="16799" />
                    <RANKING order="10" place="10" resultid="18861" />
                    <RANKING order="11" place="11" resultid="16477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9801" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19731" />
                    <RANKING order="2" place="2" resultid="19180" />
                    <RANKING order="3" place="3" resultid="17770" />
                    <RANKING order="4" place="4" resultid="18241" />
                    <RANKING order="5" place="5" resultid="18322" />
                    <RANKING order="6" place="6" resultid="19725" />
                    <RANKING order="7" place="7" resultid="17146" />
                    <RANKING order="8" place="8" resultid="18901" />
                    <RANKING order="9" place="9" resultid="18108" />
                    <RANKING order="10" place="10" resultid="17006" />
                    <RANKING order="11" place="11" resultid="16444" />
                    <RANKING order="12" place="-1" resultid="18526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9802" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18535" />
                    <RANKING order="2" place="2" resultid="18396" />
                    <RANKING order="3" place="3" resultid="17892" />
                    <RANKING order="4" place="4" resultid="19037" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19968" daytime="16:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19969" daytime="16:11" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19970" daytime="16:13" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19971" daytime="16:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19972" daytime="16:17" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19973" daytime="16:18" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19974" daytime="16:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19975" daytime="16:21" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3512" daytime="17:13" gender="M" number="18" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9832" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18197" />
                    <RANKING order="2" place="2" resultid="17296" />
                    <RANKING order="3" place="3" resultid="16601" />
                    <RANKING order="4" place="4" resultid="17301" />
                    <RANKING order="5" place="5" resultid="17875" />
                    <RANKING order="6" place="6" resultid="17289" />
                    <RANKING order="7" place="7" resultid="18716" />
                    <RANKING order="8" place="8" resultid="18257" />
                    <RANKING order="9" place="9" resultid="16641" />
                    <RANKING order="10" place="10" resultid="19310" />
                    <RANKING order="11" place="11" resultid="17500" />
                    <RANKING order="12" place="12" resultid="16618" />
                    <RANKING order="13" place="13" resultid="18435" />
                    <RANKING order="14" place="14" resultid="17956" />
                    <RANKING order="15" place="15" resultid="17283" />
                    <RANKING order="16" place="16" resultid="18248" />
                    <RANKING order="17" place="17" resultid="18664" />
                    <RANKING order="18" place="18" resultid="18313" />
                    <RANKING order="19" place="19" resultid="17951" />
                    <RANKING order="20" place="20" resultid="16940" />
                    <RANKING order="21" place="-1" resultid="17416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9833" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17869" />
                    <RANKING order="2" place="2" resultid="16742" />
                    <RANKING order="3" place="3" resultid="16704" />
                    <RANKING order="4" place="4" resultid="17529" />
                    <RANKING order="5" place="5" resultid="19748" />
                    <RANKING order="6" place="6" resultid="17119" />
                    <RANKING order="7" place="7" resultid="17588" />
                    <RANKING order="8" place="8" resultid="17483" />
                    <RANKING order="9" place="9" resultid="17155" />
                    <RANKING order="10" place="10" resultid="16858" />
                    <RANKING order="11" place="11" resultid="17248" />
                    <RANKING order="12" place="12" resultid="17961" />
                    <RANKING order="13" place="13" resultid="16783" />
                    <RANKING order="14" place="14" resultid="17983" />
                    <RANKING order="15" place="15" resultid="17362" />
                    <RANKING order="16" place="16" resultid="18179" />
                    <RANKING order="17" place="17" resultid="16925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9834" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17708" />
                    <RANKING order="2" place="2" resultid="18628" />
                    <RANKING order="3" place="3" resultid="17210" />
                    <RANKING order="4" place="4" resultid="18170" />
                    <RANKING order="5" place="5" resultid="18636" />
                    <RANKING order="6" place="6" resultid="17477" />
                    <RANKING order="7" place="7" resultid="18957" />
                    <RANKING order="8" place="8" resultid="16664" />
                    <RANKING order="9" place="9" resultid="17738" />
                    <RANKING order="10" place="10" resultid="17352" />
                    <RANKING order="11" place="11" resultid="18284" />
                    <RANKING order="12" place="12" resultid="16486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9835" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18792" />
                    <RANKING order="2" place="2" resultid="17688" />
                    <RANKING order="3" place="3" resultid="16733" />
                    <RANKING order="4" place="4" resultid="17423" />
                    <RANKING order="5" place="5" resultid="18644" />
                    <RANKING order="6" place="6" resultid="17228" />
                    <RANKING order="7" place="-1" resultid="17337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9836" agemax="20" agemin="19" name="Breedy Badger" />
                <AGEGROUP agegroupid="9837" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17494" />
                    <RANKING order="2" place="2" resultid="17262" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19994" daytime="17:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19995" daytime="17:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19996" daytime="17:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19997" daytime="17:24" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19998" daytime="17:27" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19999" daytime="17:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20000" daytime="17:33" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20001" daytime="17:36" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3545" daytime="15:12" gender="M" number="12" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9820" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17295" />
                    <RANKING order="2" place="2" resultid="18196" />
                    <RANKING order="3" place="3" resultid="19061" />
                    <RANKING order="4" place="4" resultid="17955" />
                    <RANKING order="5" place="5" resultid="16681" />
                    <RANKING order="6" place="6" resultid="18797" />
                    <RANKING order="7" place="7" resultid="18663" />
                    <RANKING order="8" place="8" resultid="17455" />
                    <RANKING order="9" place="9" resultid="18256" />
                    <RANKING order="10" place="10" resultid="17909" />
                    <RANKING order="11" place="11" resultid="18671" />
                    <RANKING order="12" place="12" resultid="18715" />
                    <RANKING order="13" place="13" resultid="17950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9821" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17430" />
                    <RANKING order="2" place="2" resultid="18619" />
                    <RANKING order="3" place="3" resultid="16672" />
                    <RANKING order="4" place="4" resultid="17603" />
                    <RANKING order="5" place="5" resultid="17751" />
                    <RANKING order="6" place="6" resultid="19127" />
                    <RANKING order="7" place="7" resultid="18912" />
                    <RANKING order="8" place="8" resultid="18142" />
                    <RANKING order="9" place="9" resultid="18187" />
                    <RANKING order="10" place="10" resultid="16711" />
                    <RANKING order="11" place="11" resultid="16782" />
                    <RANKING order="12" place="12" resultid="17369" />
                    <RANKING order="13" place="13" resultid="17154" />
                    <RANKING order="14" place="14" resultid="17903" />
                    <RANKING order="15" place="15" resultid="16426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9822" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17728" />
                    <RANKING order="2" place="2" resultid="17718" />
                    <RANKING order="3" place="3" resultid="18623" />
                    <RANKING order="4" place="4" resultid="16717" />
                    <RANKING order="5" place="5" resultid="17208" />
                    <RANKING order="6" place="6" resultid="16465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9823" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17703" />
                    <RANKING order="2" place="2" resultid="17693" />
                    <RANKING order="3" place="3" resultid="17438" />
                    <RANKING order="4" place="4" resultid="17469" />
                    <RANKING order="5" place="5" resultid="18648" />
                    <RANKING order="6" place="6" resultid="18984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9824" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17252" />
                    <RANKING order="2" place="2" resultid="19734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9825" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18612" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19911" daytime="15:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19912" daytime="15:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19913" daytime="15:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19914" daytime="15:23" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19915" daytime="15:27" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19916" daytime="15:30" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-05-08" daytime="09:30" name="Breedy Badger" number="3" warmupfrom="08:30" warmupuntil="09:20">
          <EVENTS>
            <EVENT eventid="3605" daytime="09:50" gender="M" number="21" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9895" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18198" />
                    <RANKING order="2" place="2" resultid="18717" />
                    <RANKING order="3" place="3" resultid="19063" />
                    <RANKING order="4" place="4" resultid="16642" />
                    <RANKING order="5" place="5" resultid="17876" />
                    <RANKING order="6" place="6" resultid="18258" />
                    <RANKING order="7" place="7" resultid="19311" />
                    <RANKING order="8" place="8" resultid="16602" />
                    <RANKING order="9" place="9" resultid="17302" />
                    <RANKING order="10" place="10" resultid="17290" />
                    <RANKING order="11" place="11" resultid="18673" />
                    <RANKING order="12" place="12" resultid="16619" />
                    <RANKING order="13" place="13" resultid="18436" />
                    <RANKING order="14" place="14" resultid="16682" />
                    <RANKING order="15" place="15" resultid="17541" />
                    <RANKING order="16" place="16" resultid="17284" />
                    <RANKING order="17" place="17" resultid="18207" />
                    <RANKING order="18" place="18" resultid="17910" />
                    <RANKING order="19" place="19" resultid="18314" />
                    <RANKING order="20" place="20" resultid="18665" />
                    <RANKING order="21" place="21" resultid="19103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9896" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17870" />
                    <RANKING order="2" place="2" resultid="16738" />
                    <RANKING order="3" place="3" resultid="16705" />
                    <RANKING order="4" place="4" resultid="18737" />
                    <RANKING order="5" place="5" resultid="17761" />
                    <RANKING order="6" place="6" resultid="17120" />
                    <RANKING order="7" place="7" resultid="17669" />
                    <RANKING order="8" place="8" resultid="17156" />
                    <RANKING order="9" place="9" resultid="18906" />
                    <RANKING order="10" place="10" resultid="17752" />
                    <RANKING order="11" place="11" resultid="18002" />
                    <RANKING order="12" place="12" resultid="17484" />
                    <RANKING order="13" place="13" resultid="18144" />
                    <RANKING order="14" place="14" resultid="18189" />
                    <RANKING order="15" place="15" resultid="16859" />
                    <RANKING order="16" place="16" resultid="17904" />
                    <RANKING order="17" place="17" resultid="17984" />
                    <RANKING order="18" place="18" resultid="17363" />
                    <RANKING order="19" place="19" resultid="18180" />
                    <RANKING order="20" place="20" resultid="19170" />
                    <RANKING order="21" place="21" resultid="17388" />
                    <RANKING order="22" place="-1" resultid="16784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9897" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17709" />
                    <RANKING order="2" place="2" resultid="18958" />
                    <RANKING order="3" place="3" resultid="17478" />
                    <RANKING order="4" place="4" resultid="17211" />
                    <RANKING order="5" place="5" resultid="17733" />
                    <RANKING order="6" place="6" resultid="18171" />
                    <RANKING order="7" place="7" resultid="17729" />
                    <RANKING order="8" place="8" resultid="17629" />
                    <RANKING order="9" place="9" resultid="17724" />
                    <RANKING order="10" place="10" resultid="17599" />
                    <RANKING order="11" place="11" resultid="16665" />
                    <RANKING order="12" place="12" resultid="17353" />
                    <RANKING order="13" place="13" resultid="16719" />
                    <RANKING order="14" place="14" resultid="17719" />
                    <RANKING order="15" place="15" resultid="18285" />
                    <RANKING order="16" place="16" resultid="16468" />
                    <RANKING order="17" place="17" resultid="18162" />
                    <RANKING order="18" place="18" resultid="18300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9898" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18366" />
                    <RANKING order="2" place="2" resultid="17689" />
                    <RANKING order="3" place="3" resultid="17100" />
                    <RANKING order="4" place="4" resultid="17424" />
                    <RANKING order="5" place="5" resultid="16734" />
                    <RANKING order="6" place="6" resultid="17699" />
                    <RANKING order="7" place="7" resultid="17338" />
                    <RANKING order="8" place="8" resultid="17229" />
                    <RANKING order="9" place="9" resultid="18135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9899" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9900" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19146" />
                    <RANKING order="2" place="2" resultid="17495" />
                    <RANKING order="3" place="3" resultid="16851" />
                    <RANKING order="4" place="-1" resultid="18381" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20013" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20014" daytime="09:53" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20015" daytime="09:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20016" daytime="09:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20017" daytime="09:58" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20018" daytime="10:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20019" daytime="10:01" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20020" daytime="10:03" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="20021" daytime="10:05" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="20022" daytime="10:06" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="12864" daytime="12:33" gender="M" number="27" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="EUR" value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12865" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19199" />
                    <RANKING order="2" place="2" resultid="18449" />
                    <RANKING order="3" place="3" resultid="19615" />
                    <RANKING order="4" place="4" resultid="19700" />
                    <RANKING order="5" place="5" resultid="17466" />
                    <RANKING order="6" place="6" resultid="19701" />
                    <RANKING order="7" place="7" resultid="19702" />
                    <RANKING order="8" place="8" resultid="16760" />
                    <RANKING order="9" place="9" resultid="19703" />
                    <RANKING order="10" place="10" resultid="18451" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20136" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20137" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3578" daytime="11:35" gender="M" number="25" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9901" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18199" />
                    <RANKING order="2" place="2" resultid="19064" />
                    <RANKING order="3" place="3" resultid="16620" />
                    <RANKING order="4" place="4" resultid="18437" />
                    <RANKING order="5" place="5" resultid="17297" />
                    <RANKING order="6" place="6" resultid="17291" />
                    <RANKING order="7" place="7" resultid="17285" />
                    <RANKING order="8" place="8" resultid="16643" />
                    <RANKING order="9" place="9" resultid="16603" />
                    <RANKING order="10" place="10" resultid="18259" />
                    <RANKING order="11" place="11" resultid="16683" />
                    <RANKING order="12" place="12" resultid="19228" />
                    <RANKING order="13" place="13" resultid="18446" />
                    <RANKING order="14" place="14" resultid="18250" />
                    <RANKING order="15" place="15" resultid="18674" />
                    <RANKING order="16" place="16" resultid="17501" />
                    <RANKING order="17" place="17" resultid="18718" />
                    <RANKING order="18" place="-1" resultid="17303" />
                    <RANKING order="19" place="-1" resultid="17417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9902" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18743" />
                    <RANKING order="2" place="2" resultid="16743" />
                    <RANKING order="3" place="3" resultid="16675" />
                    <RANKING order="4" place="4" resultid="17746" />
                    <RANKING order="5" place="5" resultid="17639" />
                    <RANKING order="6" place="6" resultid="16706" />
                    <RANKING order="7" place="7" resultid="17121" />
                    <RANKING order="8" place="8" resultid="17674" />
                    <RANKING order="9" place="9" resultid="17157" />
                    <RANKING order="10" place="10" resultid="16712" />
                    <RANKING order="11" place="11" resultid="17589" />
                    <RANKING order="12" place="12" resultid="16860" />
                    <RANKING order="13" place="13" resultid="17962" />
                    <RANKING order="14" place="14" resultid="17985" />
                    <RANKING order="15" place="15" resultid="17905" />
                    <RANKING order="16" place="16" resultid="17881" />
                    <RANKING order="17" place="17" resultid="17389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9903" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18172" />
                    <RANKING order="2" place="2" resultid="18428" />
                    <RANKING order="3" place="3" resultid="17965" />
                    <RANKING order="4" place="4" resultid="17734" />
                    <RANKING order="5" place="5" resultid="17742" />
                    <RANKING order="6" place="6" resultid="19269" />
                    <RANKING order="7" place="7" resultid="16666" />
                    <RANKING order="8" place="8" resultid="18286" />
                    <RANKING order="9" place="9" resultid="16720" />
                    <RANKING order="10" place="10" resultid="17609" />
                    <RANKING order="11" place="11" resultid="17193" />
                    <RANKING order="12" place="12" resultid="18959" />
                    <RANKING order="13" place="13" resultid="16469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9904" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18793" />
                    <RANKING order="2" place="2" resultid="17704" />
                    <RANKING order="3" place="3" resultid="16735" />
                    <RANKING order="4" place="4" resultid="17101" />
                    <RANKING order="5" place="5" resultid="17230" />
                    <RANKING order="6" place="6" resultid="19248" />
                    <RANKING order="7" place="7" resultid="18985" />
                    <RANKING order="8" place="8" resultid="19117" />
                    <RANKING order="9" place="9" resultid="19111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9905" agemax="20" agemin="19" name="Breedy Badger" />
                <AGEGROUP agegroupid="9906" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19100" />
                    <RANKING order="2" place="2" resultid="18383" />
                    <RANKING order="3" place="3" resultid="19094" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20051" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20052" daytime="11:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20053" daytime="11:49" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20054" daytime="11:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20055" daytime="12:01" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20056" daytime="12:07" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20057" daytime="12:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20058" daytime="12:17" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3658" daytime="10:27" gender="F" number="24" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9863" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17831" />
                    <RANKING order="2" place="2" resultid="16585" />
                    <RANKING order="3" place="3" resultid="17166" />
                    <RANKING order="4" place="4" resultid="18894" />
                    <RANKING order="5" place="5" resultid="16628" />
                    <RANKING order="6" place="6" resultid="18235" />
                    <RANKING order="7" place="7" resultid="18375" />
                    <RANKING order="8" place="8" resultid="18102" />
                    <RANKING order="9" place="9" resultid="17309" />
                    <RANKING order="10" place="10" resultid="17844" />
                    <RANKING order="11" place="11" resultid="17839" />
                    <RANKING order="12" place="12" resultid="16834" />
                    <RANKING order="13" place="13" resultid="16594" />
                    <RANKING order="14" place="14" resultid="17665" />
                    <RANKING order="15" place="15" resultid="18824" />
                    <RANKING order="16" place="16" resultid="16727" />
                    <RANKING order="17" place="17" resultid="17202" />
                    <RANKING order="18" place="18" resultid="18226" />
                    <RANKING order="19" place="19" resultid="17649" />
                    <RANKING order="20" place="20" resultid="17315" />
                    <RANKING order="21" place="21" resultid="19712" />
                    <RANKING order="22" place="22" resultid="17898" />
                    <RANKING order="23" place="23" resultid="18974" />
                    <RANKING order="24" place="24" resultid="18711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9864" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18342" />
                    <RANKING order="2" place="2" resultid="18351" />
                    <RANKING order="3" place="3" resultid="16612" />
                    <RANKING order="4" place="4" resultid="18293" />
                    <RANKING order="5" place="5" resultid="19011" />
                    <RANKING order="6" place="6" resultid="18153" />
                    <RANKING order="7" place="7" resultid="18093" />
                    <RANKING order="8" place="8" resultid="18855" />
                    <RANKING order="9" place="9" resultid="16650" />
                    <RANKING order="10" place="10" resultid="17594" />
                    <RANKING order="11" place="11" resultid="17827" />
                    <RANKING order="12" place="12" resultid="18277" />
                    <RANKING order="13" place="13" resultid="17110" />
                    <RANKING order="14" place="14" resultid="16758" />
                    <RANKING order="15" place="15" resultid="18360" />
                    <RANKING order="16" place="16" resultid="17814" />
                    <RANKING order="17" place="17" resultid="17130" />
                    <RANKING order="18" place="18" resultid="19155" />
                    <RANKING order="19" place="19" resultid="19265" />
                    <RANKING order="20" place="20" resultid="18081" />
                    <RANKING order="21" place="21" resultid="19245" />
                    <RANKING order="22" place="22" resultid="17175" />
                    <RANKING order="23" place="23" resultid="16810" />
                    <RANKING order="24" place="24" resultid="16457" />
                    <RANKING order="25" place="25" resultid="19122" />
                    <RANKING order="26" place="26" resultid="16689" />
                    <RANKING order="27" place="27" resultid="19031" />
                    <RANKING order="28" place="28" resultid="16825" />
                    <RANKING order="29" place="29" resultid="16437" />
                    <RANKING order="30" place="30" resultid="17922" />
                    <RANKING order="31" place="-1" resultid="17809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9865" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17796" />
                    <RANKING order="2" place="2" resultid="17556" />
                    <RANKING order="3" place="3" resultid="16698" />
                    <RANKING order="4" place="4" resultid="17184" />
                    <RANKING order="5" place="5" resultid="18268" />
                    <RANKING order="6" place="6" resultid="18406" />
                    <RANKING order="7" place="7" resultid="17917" />
                    <RANKING order="8" place="8" resultid="18419" />
                    <RANKING order="9" place="9" resultid="17791" />
                    <RANKING order="10" place="10" resultid="17566" />
                    <RANKING order="11" place="11" resultid="18333" />
                    <RANKING order="12" place="12" resultid="17939" />
                    <RANKING order="13" place="13" resultid="18864" />
                    <RANKING order="14" place="14" resultid="16479" />
                    <RANKING order="15" place="15" resultid="18872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9866" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17848" />
                    <RANKING order="2" place="2" resultid="17148" />
                    <RANKING order="3" place="3" resultid="18066" />
                    <RANKING order="4" place="4" resultid="16447" />
                    <RANKING order="5" place="-1" resultid="18324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9867" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18397" />
                    <RANKING order="2" place="2" resultid="17893" />
                    <RANKING order="3" place="3" resultid="16414" />
                    <RANKING order="4" place="-1" resultid="18771" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20040" daytime="10:27" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20041" daytime="10:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20042" daytime="10:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20043" daytime="10:49" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20044" daytime="10:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20045" daytime="11:01" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20046" daytime="11:07" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20047" daytime="11:13" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="20048" daytime="11:18" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="20049" daytime="11:24" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="20050" daytime="11:29" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="12862" daytime="12:22" gender="F" number="26" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="EUR" value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12863" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18452" />
                    <RANKING order="2" place="2" resultid="19704" />
                    <RANKING order="3" place="3" resultid="16762" />
                    <RANKING order="4" place="4" resultid="18454" />
                    <RANKING order="5" place="5" resultid="19202" />
                    <RANKING order="6" place="6" resultid="18456" />
                    <RANKING order="7" place="7" resultid="19705" />
                    <RANKING order="8" place="8" resultid="19706" />
                    <RANKING order="9" place="9" resultid="19203" />
                    <RANKING order="10" place="10" resultid="17233" />
                    <RANKING order="11" place="11" resultid="16489" />
                    <RANKING order="12" place="12" resultid="19707" />
                    <RANKING order="13" place="13" resultid="18836" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20134" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20135" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3617" daytime="10:08" gender="F" number="22" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9883" agemax="10" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17931" />
                    <RANKING order="2" place="2" resultid="18788" />
                    <RANKING order="3" place="3" resultid="20274" />
                    <RANKING order="4" place="4" resultid="18307" />
                    <RANKING order="5" place="5" resultid="19083" />
                    <RANKING order="6" place="6" resultid="18834" />
                    <RANKING order="7" place="7" resultid="19262" />
                    <RANKING order="8" place="8" resultid="19254" />
                    <RANKING order="9" place="9" resultid="18886" />
                    <RANKING order="10" place="10" resultid="18934" />
                    <RANKING order="11" place="11" resultid="19140" />
                    <RANKING order="12" place="12" resultid="19233" />
                    <RANKING order="13" place="13" resultid="18816" />
                    <RANKING order="14" place="14" resultid="18920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9884" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16869" />
                    <RANKING order="2" place="2" resultid="17165" />
                    <RANKING order="3" place="3" resultid="18374" />
                    <RANKING order="4" place="4" resultid="18973" />
                    <RANKING order="5" place="5" resultid="17990" />
                    <RANKING order="6" place="6" resultid="16833" />
                    <RANKING order="7" place="7" resultid="18779" />
                    <RANKING order="8" place="8" resultid="18702" />
                    <RANKING order="9" place="9" resultid="18694" />
                    <RANKING order="10" place="10" resultid="18682" />
                    <RANKING order="11" place="11" resultid="18968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9885" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19714" />
                    <RANKING order="2" place="2" resultid="18991" />
                    <RANKING order="3" place="3" resultid="17576" />
                    <RANKING order="4" place="4" resultid="17268" />
                    <RANKING order="5" place="5" resultid="17129" />
                    <RANKING order="6" place="6" resultid="19163" />
                    <RANKING order="7" place="7" resultid="17174" />
                    <RANKING order="8" place="8" resultid="19030" />
                    <RANKING order="9" place="9" resultid="16456" />
                    <RANKING order="10" place="10" resultid="16817" />
                    <RANKING order="11" place="11" resultid="16749" />
                    <RANKING order="12" place="12" resultid="17996" />
                    <RANKING order="13" place="13" resultid="18217" />
                    <RANKING order="14" place="14" resultid="17978" />
                    <RANKING order="15" place="15" resultid="18389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9886" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17916" />
                    <RANKING order="2" place="2" resultid="16636" />
                    <RANKING order="3" place="3" resultid="17561" />
                    <RANKING order="4" place="4" resultid="17943" />
                    <RANKING order="5" place="5" resultid="18054" />
                    <RANKING order="6" place="6" resultid="18405" />
                    <RANKING order="7" place="7" resultid="16844" />
                    <RANKING order="8" place="8" resultid="17183" />
                    <RANKING order="9" place="9" resultid="18418" />
                    <RANKING order="10" place="10" resultid="17781" />
                    <RANKING order="11" place="11" resultid="18128" />
                    <RANKING order="12" place="12" resultid="17346" />
                    <RANKING order="13" place="13" resultid="19197" />
                    <RANKING order="14" place="14" resultid="16877" />
                    <RANKING order="15" place="15" resultid="16802" />
                    <RANKING order="16" place="16" resultid="16478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9887" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17771" />
                    <RANKING order="2" place="2" resultid="19182" />
                    <RANKING order="3" place="3" resultid="18242" />
                    <RANKING order="4" place="4" resultid="18410" />
                    <RANKING order="5" place="5" resultid="18039" />
                    <RANKING order="6" place="6" resultid="17147" />
                    <RANKING order="7" place="7" resultid="18902" />
                    <RANKING order="8" place="8" resultid="17853" />
                    <RANKING order="9" place="9" resultid="18110" />
                    <RANKING order="10" place="10" resultid="16446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9888" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19039" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20023" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20024" daytime="10:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20025" daytime="10:11" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20026" daytime="10:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20027" daytime="10:13" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20028" daytime="10:14" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20029" daytime="10:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20030" daytime="10:16" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="20031" daytime="10:17" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3598" daytime="09:30" gender="F" number="20" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9853" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16868" />
                    <RANKING order="2" place="2" resultid="16584" />
                    <RANKING order="3" place="3" resultid="16593" />
                    <RANKING order="4" place="4" resultid="18893" />
                    <RANKING order="5" place="5" resultid="16627" />
                    <RANKING order="6" place="6" resultid="19318" />
                    <RANKING order="7" place="7" resultid="19296" />
                    <RANKING order="8" place="8" resultid="17654" />
                    <RANKING order="9" place="9" resultid="18234" />
                    <RANKING order="10" place="10" resultid="17664" />
                    <RANKING order="11" place="11" resultid="17308" />
                    <RANKING order="12" place="12" resultid="19045" />
                    <RANKING order="13" place="13" resultid="17201" />
                    <RANKING order="14" place="14" resultid="18101" />
                    <RANKING order="15" place="15" resultid="17314" />
                    <RANKING order="16" place="16" resultid="18701" />
                    <RANKING order="17" place="17" resultid="18823" />
                    <RANKING order="18" place="18" resultid="16726" />
                    <RANKING order="19" place="19" resultid="18710" />
                    <RANKING order="20" place="20" resultid="17659" />
                    <RANKING order="21" place="21" resultid="18693" />
                    <RANKING order="22" place="22" resultid="18681" />
                    <RANKING order="23" place="23" resultid="17925" />
                    <RANKING order="24" place="24" resultid="18225" />
                    <RANKING order="25" place="25" resultid="17886" />
                    <RANKING order="26" place="26" resultid="19711" />
                    <RANKING order="27" place="27" resultid="18967" />
                    <RANKING order="28" place="-1" resultid="17863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9854" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19154" />
                    <RANKING order="2" place="2" resultid="18854" />
                    <RANKING order="3" place="3" resultid="17584" />
                    <RANKING order="4" place="4" resultid="16611" />
                    <RANKING order="5" place="5" resultid="18080" />
                    <RANKING order="6" place="6" resultid="18341" />
                    <RANKING order="7" place="7" resultid="17817" />
                    <RANKING order="8" place="8" resultid="17267" />
                    <RANKING order="9" place="9" resultid="18350" />
                    <RANKING order="10" place="10" resultid="17813" />
                    <RANKING order="11" place="11" resultid="17572" />
                    <RANKING order="12" place="12" resultid="19162" />
                    <RANKING order="13" place="13" resultid="18092" />
                    <RANKING order="14" place="14" resultid="17109" />
                    <RANKING order="15" place="15" resultid="18152" />
                    <RANKING order="16" place="16" resultid="18359" />
                    <RANKING order="17" place="17" resultid="18276" />
                    <RANKING order="18" place="18" resultid="16809" />
                    <RANKING order="19" place="19" resultid="16757" />
                    <RANKING order="20" place="20" resultid="17804" />
                    <RANKING order="21" place="21" resultid="17822" />
                    <RANKING order="22" place="22" resultid="18216" />
                    <RANKING order="23" place="23" resultid="16794" />
                    <RANKING order="24" place="24" resultid="18388" />
                    <RANKING order="25" place="25" resultid="16436" />
                    <RANKING order="26" place="26" resultid="17995" />
                    <RANKING order="27" place="27" resultid="18047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9855" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16697" />
                    <RANKING order="2" place="2" resultid="18127" />
                    <RANKING order="3" place="3" resultid="18267" />
                    <RANKING order="4" place="4" resultid="16876" />
                    <RANKING order="5" place="4" resultid="18332" />
                    <RANKING order="6" place="6" resultid="19196" />
                    <RANKING order="7" place="7" resultid="17786" />
                    <RANKING order="8" place="8" resultid="16801" />
                    <RANKING order="9" place="8" resultid="17938" />
                    <RANKING order="10" place="10" resultid="18863" />
                    <RANKING order="11" place="11" resultid="18871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9856" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17776" />
                    <RANKING order="2" place="2" resultid="18409" />
                    <RANKING order="3" place="3" resultid="19181" />
                    <RANKING order="4" place="4" resultid="18323" />
                    <RANKING order="5" place="5" resultid="18109" />
                    <RANKING order="6" place="6" resultid="18065" />
                    <RANKING order="7" place="-1" resultid="16445" />
                    <RANKING order="8" place="-1" resultid="17546" />
                    <RANKING order="9" place="-1" resultid="17551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9857" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19038" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20002" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20003" daytime="09:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20004" daytime="09:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20005" daytime="09:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20006" daytime="09:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20007" daytime="09:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20008" daytime="09:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20009" daytime="09:43" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="20010" daytime="09:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="20011" daytime="09:47" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="20012" daytime="09:48" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3613" daytime="10:18" gender="M" number="23" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9925" agemax="10" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19071" />
                    <RANKING order="2" place="2" resultid="18808" />
                    <RANKING order="3" place="3" resultid="19279" />
                    <RANKING order="4" place="4" resultid="18829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9926" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18208" />
                    <RANKING order="2" place="2" resultid="19227" />
                    <RANKING order="3" place="3" resultid="18249" />
                    <RANKING order="4" place="4" resultid="18445" />
                    <RANKING order="5" place="5" resultid="17457" />
                    <RANKING order="6" place="6" resultid="18315" />
                    <RANKING order="7" place="7" resultid="18666" />
                    <RANKING order="8" place="8" resultid="19104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9927" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17624" />
                    <RANKING order="2" place="2" resultid="16674" />
                    <RANKING order="3" place="3" resultid="17432" />
                    <RANKING order="4" place="4" resultid="18738" />
                    <RANKING order="5" place="5" resultid="18907" />
                    <RANKING order="6" place="6" resultid="18914" />
                    <RANKING order="7" place="7" resultid="17604" />
                    <RANKING order="8" place="8" resultid="16785" />
                    <RANKING order="9" place="9" resultid="18190" />
                    <RANKING order="10" place="10" resultid="18145" />
                    <RANKING order="11" place="11" resultid="19089" />
                    <RANKING order="12" place="12" resultid="19129" />
                    <RANKING order="13" place="13" resultid="17364" />
                    <RANKING order="14" place="14" resultid="18181" />
                    <RANKING order="15" place="15" resultid="19171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9928" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18427" />
                    <RANKING order="2" place="2" resultid="17859" />
                    <RANKING order="3" place="3" resultid="17715" />
                    <RANKING order="4" place="4" resultid="17448" />
                    <RANKING order="5" place="5" resultid="17710" />
                    <RANKING order="6" place="6" resultid="17212" />
                    <RANKING order="7" place="7" resultid="17614" />
                    <RANKING order="8" place="8" resultid="17192" />
                    <RANKING order="9" place="9" resultid="17645" />
                    <RANKING order="10" place="10" resultid="17354" />
                    <RANKING order="11" place="11" resultid="17619" />
                    <RANKING order="12" place="12" resultid="19077" />
                    <RANKING order="13" place="13" resultid="17634" />
                    <RANKING order="14" place="14" resultid="18163" />
                    <RANKING order="15" place="15" resultid="18301" />
                    <RANKING order="16" place="16" resultid="17381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9929" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18367" />
                    <RANKING order="2" place="2" resultid="17766" />
                    <RANKING order="3" place="3" resultid="17694" />
                    <RANKING order="4" place="4" resultid="17440" />
                    <RANKING order="5" place="5" resultid="17339" />
                    <RANKING order="6" place="6" resultid="18136" />
                    <RANKING order="7" place="7" resultid="19116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9930" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17409" />
                    <RANKING order="2" place="2" resultid="17679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9931" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19051" />
                    <RANKING order="2" place="2" resultid="19135" />
                    <RANKING order="3" place="3" resultid="19189" />
                    <RANKING order="4" place="4" resultid="18951" />
                    <RANKING order="5" place="5" resultid="17496" />
                    <RANKING order="6" place="6" resultid="16852" />
                    <RANKING order="7" place="7" resultid="18945" />
                    <RANKING order="8" place="8" resultid="17328" />
                    <RANKING order="9" place="-1" resultid="19258" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20032" daytime="10:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20033" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20034" daytime="10:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20035" daytime="10:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20036" daytime="10:23" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20037" daytime="10:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20038" daytime="10:24" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20039" daytime="10:25" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-05-08" daytime="13:30" name="Breedy Badger" number="4">
          <EVENTS>
            <EVENT eventid="3530" daytime="14:34" gender="M" number="33" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9913" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19066" />
                    <RANKING order="2" place="2" resultid="18201" />
                    <RANKING order="3" place="3" resultid="16621" />
                    <RANKING order="4" place="4" resultid="18676" />
                    <RANKING order="5" place="5" resultid="17292" />
                    <RANKING order="6" place="6" resultid="16644" />
                    <RANKING order="7" place="7" resultid="17542" />
                    <RANKING order="8" place="8" resultid="18439" />
                    <RANKING order="9" place="9" resultid="16604" />
                    <RANKING order="10" place="10" resultid="16684" />
                    <RANKING order="11" place="11" resultid="17538" />
                    <RANKING order="12" place="12" resultid="18261" />
                    <RANKING order="13" place="13" resultid="17286" />
                    <RANKING order="14" place="14" resultid="17304" />
                    <RANKING order="15" place="15" resultid="19229" />
                    <RANKING order="16" place="16" resultid="18252" />
                    <RANKING order="17" place="17" resultid="18448" />
                    <RANKING order="18" place="18" resultid="17502" />
                    <RANKING order="19" place="19" resultid="17877" />
                    <RANKING order="20" place="20" resultid="18210" />
                    <RANKING order="21" place="21" resultid="19312" />
                    <RANKING order="22" place="22" resultid="17911" />
                    <RANKING order="23" place="23" resultid="18317" />
                    <RANKING order="24" place="24" resultid="17459" />
                    <RANKING order="25" place="25" resultid="18668" />
                    <RANKING order="26" place="26" resultid="17419" />
                    <RANKING order="27" place="27" resultid="19303" />
                    <RANKING order="28" place="28" resultid="19106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9914" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18745" />
                    <RANKING order="2" place="2" resultid="19282" />
                    <RANKING order="3" place="3" resultid="18740" />
                    <RANKING order="4" place="4" resultid="17748" />
                    <RANKING order="5" place="5" resultid="17434" />
                    <RANKING order="6" place="6" resultid="17123" />
                    <RANKING order="7" place="7" resultid="17757" />
                    <RANKING order="8" place="8" resultid="17530" />
                    <RANKING order="9" place="9" resultid="17753" />
                    <RANKING order="10" place="10" resultid="19287" />
                    <RANKING order="11" place="11" resultid="17159" />
                    <RANKING order="12" place="12" resultid="18147" />
                    <RANKING order="13" place="13" resultid="17906" />
                    <RANKING order="14" place="14" resultid="16787" />
                    <RANKING order="15" place="15" resultid="18003" />
                    <RANKING order="16" place="16" resultid="18192" />
                    <RANKING order="17" place="17" resultid="18916" />
                    <RANKING order="18" place="18" resultid="17486" />
                    <RANKING order="19" place="19" resultid="17963" />
                    <RANKING order="20" place="20" resultid="19131" />
                    <RANKING order="21" place="21" resultid="17371" />
                    <RANKING order="22" place="22" resultid="16861" />
                    <RANKING order="23" place="23" resultid="17365" />
                    <RANKING order="24" place="24" resultid="19090" />
                    <RANKING order="25" place="25" resultid="18183" />
                    <RANKING order="26" place="26" resultid="19173" />
                    <RANKING order="27" place="27" resultid="17391" />
                    <RANKING order="28" place="-1" resultid="17625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9915" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18430" />
                    <RANKING order="2" place="2" resultid="17479" />
                    <RANKING order="3" place="3" resultid="17735" />
                    <RANKING order="4" place="4" resultid="17615" />
                    <RANKING order="5" place="5" resultid="17630" />
                    <RANKING order="6" place="6" resultid="17213" />
                    <RANKING order="7" place="7" resultid="17356" />
                    <RANKING order="8" place="8" resultid="17451" />
                    <RANKING order="9" place="9" resultid="16668" />
                    <RANKING order="10" place="10" resultid="19079" />
                    <RANKING order="11" place="11" resultid="16470" />
                    <RANKING order="12" place="12" resultid="17195" />
                    <RANKING order="13" place="13" resultid="17635" />
                    <RANKING order="14" place="14" resultid="18287" />
                    <RANKING order="15" place="15" resultid="18165" />
                    <RANKING order="16" place="16" resultid="17383" />
                    <RANKING order="17" place="17" resultid="18303" />
                    <RANKING order="18" place="-1" resultid="18960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9916" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18368" />
                    <RANKING order="2" place="2" resultid="19240" />
                    <RANKING order="3" place="3" resultid="17472" />
                    <RANKING order="4" place="4" resultid="17767" />
                    <RANKING order="5" place="5" resultid="17426" />
                    <RANKING order="6" place="6" resultid="17442" />
                    <RANKING order="7" place="7" resultid="19112" />
                    <RANKING order="8" place="8" resultid="19250" />
                    <RANKING order="9" place="9" resultid="17340" />
                    <RANKING order="10" place="10" resultid="17232" />
                    <RANKING order="11" place="11" resultid="19118" />
                    <RANKING order="12" place="12" resultid="18138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9917" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17411" />
                    <RANKING order="2" place="2" resultid="17680" />
                    <RANKING order="3" place="3" resultid="17685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9918" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19052" />
                    <RANKING order="2" place="2" resultid="19136" />
                    <RANKING order="3" place="3" resultid="19101" />
                    <RANKING order="4" place="4" resultid="16853" />
                    <RANKING order="5" place="5" resultid="18952" />
                    <RANKING order="6" place="6" resultid="18946" />
                    <RANKING order="7" place="7" resultid="19191" />
                    <RANKING order="8" place="8" resultid="19095" />
                    <RANKING order="9" place="9" resultid="17330" />
                    <RANKING order="10" place="10" resultid="18941" />
                    <RANKING order="11" place="-1" resultid="18382" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20100" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20101" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20102" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20103" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20104" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20105" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20106" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20107" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="20108" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="20109" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="20110" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="20111" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="20112" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3523" daytime="14:10" gender="F" number="32" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9873" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17510" />
                    <RANKING order="2" place="2" resultid="16586" />
                    <RANKING order="3" place="3" resultid="17836" />
                    <RANKING order="4" place="4" resultid="18895" />
                    <RANKING order="5" place="5" resultid="19046" />
                    <RANKING order="6" place="6" resultid="19319" />
                    <RANKING order="7" place="7" resultid="16629" />
                    <RANKING order="8" place="8" resultid="16595" />
                    <RANKING order="9" place="9" resultid="17168" />
                    <RANKING order="10" place="10" resultid="17310" />
                    <RANKING order="11" place="11" resultid="17840" />
                    <RANKING order="12" place="12" resultid="18103" />
                    <RANKING order="13" place="13" resultid="19297" />
                    <RANKING order="14" place="14" resultid="18377" />
                    <RANKING order="15" place="15" resultid="18237" />
                    <RANKING order="16" place="16" resultid="17204" />
                    <RANKING order="17" place="17" resultid="16728" />
                    <RANKING order="18" place="18" resultid="18826" />
                    <RANKING order="19" place="19" resultid="17316" />
                    <RANKING order="20" place="20" resultid="17506" />
                    <RANKING order="21" place="21" resultid="17514" />
                    <RANKING order="22" place="22" resultid="18228" />
                    <RANKING order="23" place="23" resultid="18712" />
                    <RANKING order="24" place="24" resultid="18975" />
                    <RANKING order="25" place="25" resultid="18781" />
                    <RANKING order="26" place="26" resultid="17650" />
                    <RANKING order="27" place="27" resultid="19713" />
                    <RANKING order="28" place="28" resultid="17927" />
                    <RANKING order="29" place="29" resultid="18704" />
                    <RANKING order="30" place="30" resultid="17887" />
                    <RANKING order="31" place="31" resultid="18696" />
                    <RANKING order="32" place="32" resultid="18969" />
                    <RANKING order="33" place="33" resultid="18684" />
                    <RANKING order="34" place="34" resultid="19291" />
                    <RANKING order="35" place="35" resultid="17864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9874" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16613" />
                    <RANKING order="2" place="2" resultid="18343" />
                    <RANKING order="3" place="3" resultid="18352" />
                    <RANKING order="4" place="4" resultid="18856" />
                    <RANKING order="5" place="5" resultid="19299" />
                    <RANKING order="6" place="6" resultid="18295" />
                    <RANKING order="7" place="7" resultid="17585" />
                    <RANKING order="8" place="8" resultid="17577" />
                    <RANKING order="9" place="9" resultid="17269" />
                    <RANKING order="10" place="10" resultid="19012" />
                    <RANKING order="11" place="11" resultid="18278" />
                    <RANKING order="12" place="12" resultid="17828" />
                    <RANKING order="13" place="13" resultid="18095" />
                    <RANKING order="14" place="14" resultid="18993" />
                    <RANKING order="15" place="15" resultid="18361" />
                    <RANKING order="16" place="16" resultid="17595" />
                    <RANKING order="17" place="17" resultid="16759" />
                    <RANKING order="18" place="18" resultid="18155" />
                    <RANKING order="19" place="19" resultid="16811" />
                    <RANKING order="20" place="20" resultid="19267" />
                    <RANKING order="21" place="21" resultid="18082" />
                    <RANKING order="22" place="22" resultid="17132" />
                    <RANKING order="23" place="23" resultid="19164" />
                    <RANKING order="24" place="24" resultid="16796" />
                    <RANKING order="25" place="25" resultid="17112" />
                    <RANKING order="26" place="26" resultid="19123" />
                    <RANKING order="27" place="27" resultid="19246" />
                    <RANKING order="28" place="28" resultid="17805" />
                    <RANKING order="29" place="29" resultid="17177" />
                    <RANKING order="30" place="30" resultid="16691" />
                    <RANKING order="31" place="31" resultid="18390" />
                    <RANKING order="32" place="32" resultid="16439" />
                    <RANKING order="33" place="33" resultid="17823" />
                    <RANKING order="34" place="34" resultid="16827" />
                    <RANKING order="35" place="35" resultid="16819" />
                    <RANKING order="36" place="36" resultid="16751" />
                    <RANKING order="37" place="37" resultid="18219" />
                    <RANKING order="38" place="38" resultid="17997" />
                    <RANKING order="39" place="39" resultid="18048" />
                    <RANKING order="40" place="40" resultid="17979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9875" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17186" />
                    <RANKING order="2" place="2" resultid="17562" />
                    <RANKING order="3" place="3" resultid="16637" />
                    <RANKING order="4" place="4" resultid="17944" />
                    <RANKING order="5" place="5" resultid="16699" />
                    <RANKING order="6" place="6" resultid="17782" />
                    <RANKING order="7" place="7" resultid="18270" />
                    <RANKING order="8" place="8" resultid="18129" />
                    <RANKING order="9" place="9" resultid="16845" />
                    <RANKING order="10" place="10" resultid="17347" />
                    <RANKING order="11" place="11" resultid="17792" />
                    <RANKING order="12" place="12" resultid="18056" />
                    <RANKING order="13" place="13" resultid="18074" />
                    <RANKING order="14" place="14" resultid="19198" />
                    <RANKING order="15" place="15" resultid="18334" />
                    <RANKING order="16" place="16" resultid="17567" />
                    <RANKING order="17" place="17" resultid="18865" />
                    <RANKING order="18" place="18" resultid="16803" />
                    <RANKING order="19" place="19" resultid="16878" />
                    <RANKING order="20" place="20" resultid="18873" />
                    <RANKING order="21" place="21" resultid="16481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9876" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18243" />
                    <RANKING order="2" place="2" resultid="17552" />
                    <RANKING order="3" place="3" resultid="19184" />
                    <RANKING order="4" place="4" resultid="18904" />
                    <RANKING order="5" place="5" resultid="17772" />
                    <RANKING order="6" place="6" resultid="17150" />
                    <RANKING order="7" place="7" resultid="18041" />
                    <RANKING order="8" place="8" resultid="17854" />
                    <RANKING order="9" place="9" resultid="18112" />
                    <RANKING order="10" place="10" resultid="18067" />
                    <RANKING order="11" place="11" resultid="16449" />
                    <RANKING order="12" place="-1" resultid="17547" />
                    <RANKING order="13" place="-1" resultid="18326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9877" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19040" />
                    <RANKING order="2" place="2" resultid="16417" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20085" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20086" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20087" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20088" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20089" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20090" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20091" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20092" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="20093" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="20094" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="20095" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="20096" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="20097" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="20098" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="20099" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3519" daytime="13:59" gender="M" number="31" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9932" agemax="10" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19280" />
                    <RANKING order="2" place="2" resultid="19072" />
                    <RANKING order="3" place="3" resultid="18809" />
                    <RANKING order="4" place="4" resultid="17463" />
                    <RANKING order="5" place="5" resultid="18830" />
                    <RANKING order="6" place="6" resultid="17489" />
                    <RANKING order="7" place="7" resultid="19306" />
                    <RANKING order="8" place="8" resultid="17974" />
                    <RANKING order="9" place="-1" resultid="17970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9933" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17957" />
                    <RANKING order="2" place="2" resultid="19065" />
                    <RANKING order="3" place="3" resultid="18200" />
                    <RANKING order="4" place="4" resultid="17298" />
                    <RANKING order="5" place="5" resultid="17458" />
                    <RANKING order="6" place="6" resultid="18667" />
                    <RANKING order="7" place="7" resultid="18675" />
                    <RANKING order="8" place="8" resultid="18260" />
                    <RANKING order="9" place="9" resultid="18438" />
                    <RANKING order="10" place="10" resultid="18251" />
                    <RANKING order="11" place="11" resultid="19105" />
                    <RANKING order="12" place="12" resultid="18316" />
                    <RANKING order="13" place="13" resultid="18447" />
                    <RANKING order="14" place="14" resultid="17418" />
                    <RANKING order="15" place="15" resultid="18209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9934" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17534" />
                    <RANKING order="2" place="2" resultid="17433" />
                    <RANKING order="3" place="3" resultid="17605" />
                    <RANKING order="4" place="4" resultid="16676" />
                    <RANKING order="5" place="5" resultid="17485" />
                    <RANKING order="6" place="6" resultid="18191" />
                    <RANKING order="7" place="7" resultid="18739" />
                    <RANKING order="8" place="8" resultid="18915" />
                    <RANKING order="9" place="9" resultid="17370" />
                    <RANKING order="10" place="10" resultid="18146" />
                    <RANKING order="11" place="11" resultid="19130" />
                    <RANKING order="12" place="12" resultid="17122" />
                    <RANKING order="13" place="13" resultid="17158" />
                    <RANKING order="14" place="14" resultid="16713" />
                    <RANKING order="15" place="15" resultid="19172" />
                    <RANKING order="16" place="16" resultid="16786" />
                    <RANKING order="17" place="17" resultid="18182" />
                    <RANKING order="18" place="18" resultid="17390" />
                    <RANKING order="19" place="19" resultid="17882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9935" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18173" />
                    <RANKING order="2" place="2" resultid="19078" />
                    <RANKING order="3" place="3" resultid="17450" />
                    <RANKING order="4" place="4" resultid="18280" />
                    <RANKING order="5" place="5" resultid="17355" />
                    <RANKING order="6" place="6" resultid="17382" />
                    <RANKING order="7" place="7" resultid="18302" />
                    <RANKING order="8" place="8" resultid="18164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9936" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17695" />
                    <RANKING order="2" place="2" resultid="17441" />
                    <RANKING order="3" place="3" resultid="19249" />
                    <RANKING order="4" place="4" resultid="17690" />
                    <RANKING order="5" place="5" resultid="18986" />
                    <RANKING order="6" place="6" resultid="17471" />
                    <RANKING order="7" place="7" resultid="17425" />
                    <RANKING order="8" place="8" resultid="18137" />
                    <RANKING order="9" place="9" resultid="17231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9937" agemax="20" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9938" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19190" />
                    <RANKING order="2" place="2" resultid="17114" />
                    <RANKING order="3" place="3" resultid="18940" />
                    <RANKING order="4" place="4" resultid="17329" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20076" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20077" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20078" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20079" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20080" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20081" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20082" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20083" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="20084" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3514" daytime="13:48" gender="F" number="30" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9889" agemax="10" agemin="-1" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18789" />
                    <RANKING order="2" place="2" resultid="19263" />
                    <RANKING order="3" place="3" resultid="17932" />
                    <RANKING order="4" place="4" resultid="19141" />
                    <RANKING order="5" place="5" resultid="18887" />
                    <RANKING order="6" place="6" resultid="18308" />
                    <RANKING order="7" place="7" resultid="19084" />
                    <RANKING order="8" place="8" resultid="18784" />
                    <RANKING order="9" place="9" resultid="19255" />
                    <RANKING order="10" place="10" resultid="19222" />
                    <RANKING order="11" place="11" resultid="19177" />
                    <RANKING order="12" place="12" resultid="19234" />
                    <RANKING order="13" place="13" resultid="18921" />
                    <RANKING order="14" place="14" resultid="18935" />
                    <RANKING order="15" place="15" resultid="18835" />
                    <RANKING order="16" place="16" resultid="18817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9890" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16836" />
                    <RANKING order="2" place="2" resultid="17899" />
                    <RANKING order="3" place="3" resultid="18703" />
                    <RANKING order="4" place="4" resultid="17203" />
                    <RANKING order="5" place="5" resultid="18780" />
                    <RANKING order="6" place="6" resultid="17518" />
                    <RANKING order="7" place="7" resultid="18236" />
                    <RANKING order="8" place="8" resultid="18695" />
                    <RANKING order="9" place="9" resultid="17526" />
                    <RANKING order="10" place="10" resultid="17926" />
                    <RANKING order="11" place="11" resultid="18227" />
                    <RANKING order="12" place="12" resultid="18376" />
                    <RANKING order="13" place="13" resultid="18683" />
                    <RANKING order="14" place="14" resultid="18962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9891" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19266" />
                    <RANKING order="2" place="2" resultid="18294" />
                    <RANKING order="3" place="3" resultid="16795" />
                    <RANKING order="4" place="4" resultid="16651" />
                    <RANKING order="5" place="5" resultid="17176" />
                    <RANKING order="6" place="6" resultid="17131" />
                    <RANKING order="7" place="7" resultid="16818" />
                    <RANKING order="8" place="8" resultid="18154" />
                    <RANKING order="9" place="9" resultid="16690" />
                    <RANKING order="10" place="10" resultid="16438" />
                    <RANKING order="11" place="11" resultid="19032" />
                    <RANKING order="12" place="12" resultid="16459" />
                    <RANKING order="13" place="13" resultid="17111" />
                    <RANKING order="14" place="14" resultid="16826" />
                    <RANKING order="15" place="15" resultid="18218" />
                    <RANKING order="16" place="16" resultid="17923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9892" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17918" />
                    <RANKING order="2" place="2" resultid="18407" />
                    <RANKING order="3" place="3" resultid="18055" />
                    <RANKING order="4" place="4" resultid="17185" />
                    <RANKING order="5" place="5" resultid="18073" />
                    <RANKING order="6" place="6" resultid="18269" />
                    <RANKING order="7" place="7" resultid="16480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9893" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18412" />
                    <RANKING order="2" place="2" resultid="17149" />
                    <RANKING order="3" place="3" resultid="18111" />
                    <RANKING order="4" place="4" resultid="18040" />
                    <RANKING order="5" place="5" resultid="17849" />
                    <RANKING order="6" place="6" resultid="16448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9894" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16416" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20068" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20069" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20070" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20071" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="20072" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="20073" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="20074" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="20075" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1081" daytime="15:16" gender="M" number="35" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9919" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9920" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16744" />
                    <RANKING order="2" place="2" resultid="17762" />
                    <RANKING order="3" place="3" resultid="16677" />
                    <RANKING order="4" place="4" resultid="18741" />
                    <RANKING order="5" place="5" resultid="16701" />
                    <RANKING order="6" place="6" resultid="17522" />
                    <RANKING order="7" place="7" resultid="16708" />
                    <RANKING order="8" place="8" resultid="17675" />
                    <RANKING order="9" place="9" resultid="17670" />
                    <RANKING order="10" place="10" resultid="17590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9921" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17966" />
                    <RANKING order="2" place="2" resultid="17730" />
                    <RANKING order="3" place="3" resultid="18174" />
                    <RANKING order="4" place="4" resultid="17214" />
                    <RANKING order="5" place="5" resultid="17743" />
                    <RANKING order="6" place="6" resultid="16721" />
                    <RANKING order="7" place="7" resultid="17600" />
                    <RANKING order="8" place="8" resultid="16471" />
                    <RANKING order="9" place="-1" resultid="17739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9922" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17705" />
                    <RANKING order="2" place="2" resultid="18794" />
                    <RANKING order="3" place="3" resultid="16736" />
                    <RANKING order="4" place="4" resultid="17103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9923" agemax="20" agemin="19" name="Breedy Badger" />
                <AGEGROUP agegroupid="9924" agemax="-1" agemin="21" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19147" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20116" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20117" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20118" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="20119" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3636" daytime="14:55" gender="F" number="34" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9878" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17832" />
                    <RANKING order="2" place="2" resultid="17655" />
                    <RANKING order="3" place="3" resultid="17660" />
                    <RANKING order="4" place="4" resultid="16837" />
                    <RANKING order="5" place="5" resultid="18825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9879" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18344" />
                    <RANKING order="2" place="2" resultid="18353" />
                    <RANKING order="3" place="3" resultid="17270" />
                    <RANKING order="4" place="4" resultid="19156" />
                    <RANKING order="5" place="5" resultid="16646" />
                    <RANKING order="6" place="6" resultid="16460" />
                    <RANKING order="7" place="7" resultid="19033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9880" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17946" />
                    <RANKING order="2" place="2" resultid="18421" />
                    <RANKING order="3" place="3" resultid="18335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9881" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9882" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18399" />
                    <RANKING order="2" place="2" resultid="16418" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20113" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20114" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20115" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3586" daytime="13:30" gender="F" number="28" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9868" agemax="12" agemin="11" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16870" />
                    <RANKING order="2" place="2" resultid="17167" />
                    <RANKING order="3" place="3" resultid="17991" />
                    <RANKING order="4" place="4" resultid="16835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9869" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17818" />
                    <RANKING order="2" place="2" resultid="18992" />
                    <RANKING order="3" place="3" resultid="17801" />
                    <RANKING order="4" place="4" resultid="16750" />
                    <RANKING order="5" place="5" resultid="18094" />
                    <RANKING order="6" place="6" resultid="16458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9870" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17797" />
                    <RANKING order="2" place="2" resultid="16631" />
                    <RANKING order="3" place="3" resultid="17557" />
                    <RANKING order="4" place="4" resultid="17787" />
                    <RANKING order="5" place="-1" resultid="18420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9871" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19285" />
                    <RANKING order="2" place="2" resultid="19183" />
                    <RANKING order="3" place="3" resultid="18903" />
                    <RANKING order="4" place="-1" resultid="18325" />
                    <RANKING order="5" place="-1" resultid="18411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9872" agemax="-1" agemin="19" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18398" />
                    <RANKING order="2" place="-1" resultid="16415" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20063" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20064" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="20065" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3588" daytime="13:41" gender="M" number="29" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9907" agemax="12" agemin="11" name="Breedy Badger" />
                <AGEGROUP agegroupid="9908" agemax="14" agemin="13" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18744" />
                    <RANKING order="2" place="2" resultid="17640" />
                    <RANKING order="3" place="3" resultid="17747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9909" agemax="16" agemin="15" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17725" />
                    <RANKING order="2" place="2" resultid="16667" />
                    <RANKING order="3" place="3" resultid="17610" />
                    <RANKING order="4" place="4" resultid="18429" />
                    <RANKING order="5" place="5" resultid="17449" />
                    <RANKING order="6" place="6" resultid="17720" />
                    <RANKING order="7" place="7" resultid="17620" />
                    <RANKING order="8" place="8" resultid="17194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9910" agemax="18" agemin="17" name="Breedy Badger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17102" />
                    <RANKING order="2" place="2" resultid="17700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9911" agemax="20" agemin="19" name="Breedy Badger" />
                <AGEGROUP agegroupid="9912" agemax="-1" agemin="21" name="Breedy Badger" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="20066" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="20067" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="TTCI" nation="AUT" region="TLSV" clubid="18747" swrid="89752" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" athleteid="18764">
              <RESULTS>
                <RESULT eventid="3547" points="125" swimtime="00:00:54.01" resultid="18765" heatid="19835" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="3570" points="105" swimtime="00:03:59.05" resultid="18766" heatid="19874" lane="4" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" athleteid="18770">
              <RESULTS>
                <RESULT comment=" - Start vor dem Startsignal (Zeit: 11:02)" eventid="3658" status="DSQ" swimtime="00:06:14.47" resultid="18771" heatid="20042" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="200" swimtime="00:02:54.94" />
                    <SPLIT distance="300" swimtime="00:04:35.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="4703559" athleteid="18772">
              <RESULTS>
                <RESULT comment=" - Start vor dem Startsignal (Zeit: 14:06)" eventid="3649" status="DSQ" swimtime="00:02:46.14" resultid="18773" heatid="19893" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="303" swimtime="00:00:31.11" resultid="18774" heatid="19953" lane="8" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" athleteid="18750">
              <RESULTS>
                <RESULT eventid="3570" points="167" reactiontime="+71" swimtime="00:03:24.81" resultid="18751" heatid="19878" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="197" swimtime="00:00:40.77" resultid="18752" heatid="19925" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" athleteid="18756">
              <RESULTS>
                <RESULT eventid="3570" points="221" reactiontime="+81" swimtime="00:03:06.62" resultid="18757" heatid="19878" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="280" swimtime="00:00:36.23" resultid="18758" heatid="19925" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" athleteid="18753">
              <RESULTS>
                <RESULT eventid="3570" points="198" swimtime="00:03:13.72" resultid="18754" heatid="19878" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="261" swimtime="00:00:37.12" resultid="18755" heatid="19925" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BZN" nation="ITA" clubid="18460" swrid="82616" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2001-07-09" firstname="Julia4" gender="M" lastname="Janke-Frosch4" nation="ITA" swrid="4841381" athleteid="18613">
              <RESULTS>
                <RESULT eventid="3551" points="536" swimtime="00:00:29.58" resultid="18614" heatid="19852" lane="7" entrytime="00:00:29.01" />
                <RESULT eventid="3649" points="482" reactiontime="+52" swimtime="00:02:10.09" resultid="18615" heatid="19896" lane="4" entrytime="00:02:11.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="484" swimtime="00:00:26.63" resultid="18616" heatid="19958" lane="1" entrytime="00:00:26.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-07-26" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4823062" athleteid="18541">
              <RESULTS>
                <RESULT eventid="3639" points="406" swimtime="00:02:50.26" resultid="18542" heatid="19817" lane="4" entrytime="00:02:48.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="422" reactiontime="+54" swimtime="00:02:30.56" resultid="18543" heatid="19883" lane="1" entrytime="00:02:30.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="446" swimtime="00:00:31.05" resultid="18544" heatid="19931" lane="8" entrytime="00:00:31.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-05-10" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4707999" athleteid="18505">
              <RESULTS>
                <RESULT eventid="3621" points="422" reactiontime="+77" swimtime="00:01:25.89" resultid="18506" heatid="19861" lane="6" entrytime="00:01:23.15" />
                <RESULT eventid="3555" points="362" reactiontime="+64" swimtime="00:01:18.61" resultid="18507" heatid="19973" lane="8" entrytime="00:01:14.39" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-05-15" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4517242" athleteid="18523">
              <RESULTS>
                <RESULT eventid="3639" points="646" reactiontime="+55" swimtime="00:02:25.91" resultid="18524" heatid="19822" lane="3" entrytime="00:02:22.52">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="627" swimtime="00:00:31.60" resultid="18525" heatid="19844" lane="4" entrytime="00:00:30.40" />
                <RESULT eventid="3555" status="DNS" swimtime="00:00:00.00" resultid="18526" heatid="19975" lane="5" entrytime="00:01:04.00" />
                <RESULT eventid="3505" points="548" swimtime="00:02:32.50" resultid="18527" heatid="19993" lane="3" entrytime="00:02:22.32">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="657" swimtime="00:00:27.29" resultid="18657" heatid="19937" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="15921" points="609" swimtime="00:00:27.99" resultid="20151" heatid="20120" lane="4" late="yes" />
                <RESULT eventid="15972" points="577" swimtime="00:00:28.49" resultid="20152" heatid="20122" lane="4" late="yes" />
                <RESULT eventid="15975" points="580" swimtime="00:00:28.45" resultid="20153" heatid="20124" lane="4" late="yes" />
                <RESULT eventid="15978" points="600" swimtime="00:00:28.13" resultid="20155" heatid="20126" lane="4" late="yes" />
                <RESULT eventid="15981" points="622" swimtime="00:00:27.79" resultid="20156" heatid="20128" lane="4" late="yes" />
                <RESULT eventid="15984" points="669" swimtime="00:00:27.12" resultid="20157" heatid="20130" lane="4" late="yes" />
                <RESULT eventid="15987" points="653" swimtime="00:00:27.35" resultid="20158" heatid="20132" lane="4" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-11-08" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4199604" athleteid="18590">
              <RESULTS>
                <RESULT eventid="3639" points="483" reactiontime="+73" swimtime="00:02:40.78" resultid="18591" heatid="19821" lane="1" entrytime="00:02:36.66">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="494" reactiontime="+76" swimtime="00:01:21.51" resultid="18592" heatid="19863" lane="8" entrytime="00:01:18.97" />
                <RESULT eventid="3538" points="488" reactiontime="+61" swimtime="00:02:57.95" resultid="18593" heatid="19910" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-11-03" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4712835" athleteid="18641">
              <RESULTS>
                <RESULT eventid="3551" points="401" swimtime="00:00:32.59" resultid="18642" heatid="19850" lane="4" entrytime="00:00:31.89" />
                <RESULT eventid="3594" points="420" swimtime="00:00:27.91" resultid="18643" heatid="19955" lane="3" entrytime="00:00:27.56" />
                <RESULT eventid="3512" points="386" swimtime="00:02:33.70" resultid="18644" heatid="20001" lane="8" entrytime="00:02:21.13">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-06" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4650018" athleteid="18557">
              <RESULTS>
                <RESULT eventid="3570" points="439" reactiontime="+84" swimtime="00:02:28.55" resultid="18558" heatid="19883" lane="6" entrytime="00:02:28.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="419" swimtime="00:00:31.70" resultid="18559" heatid="19930" lane="4" entrytime="00:00:31.40" />
                <RESULT eventid="3555" points="432" swimtime="00:01:14.12" resultid="18560" heatid="19973" lane="1" entrytime="00:01:13.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-21" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4823064" athleteid="18617">
              <RESULTS>
                <RESULT eventid="3628" points="431" swimtime="00:01:17.55" resultid="18618" heatid="19870" lane="4" entrytime="00:01:19.56" />
                <RESULT eventid="3545" points="437" swimtime="00:02:47.65" resultid="18619" heatid="19915" lane="3" entrytime="00:02:46.65">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="263" swimtime="00:00:32.61" resultid="18620" heatid="19951" lane="1" entrytime="00:00:32.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-09-08" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5089280" athleteid="18497">
              <RESULTS>
                <RESULT eventid="3621" points="301" reactiontime="+74" swimtime="00:01:36.14" resultid="18498" heatid="19856" lane="1" entrytime="00:01:41.11" />
                <RESULT eventid="3570" points="310" reactiontime="+67" swimtime="00:02:46.79" resultid="18499" heatid="19877" lane="7" entrytime="00:02:58.78">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="319" swimtime="00:00:34.71" resultid="18500" heatid="19924" lane="8" entrytime="00:00:36.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-02-11" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4316130" athleteid="18609">
              <RESULTS>
                <RESULT eventid="9711" points="485" reactiontime="+73" swimtime="00:02:25.07" resultid="18610" heatid="19832" lane="6" entrytime="00:02:13.35">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="597" reactiontime="+57" swimtime="00:01:09.57" resultid="18611" heatid="19872" lane="4" entrytime="00:01:02.65" />
                <RESULT eventid="3545" points="561" reactiontime="+61" swimtime="00:02:34.29" resultid="18612" heatid="19916" lane="4" entrytime="00:02:14.14">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-03-28" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4649989" athleteid="18573">
              <RESULTS>
                <RESULT eventid="3639" points="519" reactiontime="+76" swimtime="00:02:36.89" resultid="18574" heatid="19822" lane="1" entrytime="00:02:33.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="506" reactiontime="+75" swimtime="00:02:21.69" resultid="18575" heatid="19887" lane="6" entrytime="00:02:15.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="468" swimtime="00:01:12.20" resultid="18576" heatid="19973" lane="5" entrytime="00:01:11.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-09-15" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4426767" athleteid="18565">
              <RESULTS>
                <RESULT eventid="3621" points="485" reactiontime="+71" swimtime="00:01:22.01" resultid="18566" heatid="19862" lane="1" entrytime="00:01:21.00" />
                <RESULT eventid="3538" points="464" reactiontime="+92" swimtime="00:03:00.95" resultid="18567" heatid="19910" lane="8" entrytime="00:02:50.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="466" swimtime="00:00:30.60" resultid="18568" heatid="19933" lane="1" entrytime="00:00:30.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-08-08" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4708015" athleteid="18545">
              <RESULTS>
                <RESULT eventid="3547" points="350" swimtime="00:00:38.39" resultid="18546" heatid="19841" lane="4" entrytime="00:00:36.60" />
                <RESULT eventid="3570" points="360" swimtime="00:02:38.70" resultid="18547" heatid="19883" lane="3" entrytime="00:02:28.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="399" swimtime="00:00:32.21" resultid="18548" heatid="19930" lane="7" entrytime="00:00:31.52" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-03-16" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4938258" athleteid="18629">
              <RESULTS>
                <RESULT eventid="3551" points="321" swimtime="00:00:35.11" resultid="18630" heatid="19849" lane="4" entrytime="00:00:34.56" />
                <RESULT comment=" - Aktiver Delphinbeinschlag (Zeit: 12:44)" eventid="3628" reactiontime="+71" status="DSQ" swimtime="00:01:25.76" resultid="18631" heatid="19869" lane="6" entrytime="00:01:22.24" />
                <RESULT eventid="3594" points="348" swimtime="00:00:29.71" resultid="18632" heatid="19952" lane="5" entrytime="00:00:29.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-06-14" firstname="Julia2" gender="M" lastname="Janke-Frosch2" nation="ITA" swrid="4900639" athleteid="18621">
              <RESULTS>
                <RESULT eventid="3628" points="459" reactiontime="+50" swimtime="00:01:15.89" resultid="18622" heatid="19871" lane="3" entrytime="00:01:15.01" />
                <RESULT eventid="3545" points="445" reactiontime="+53" swimtime="00:02:46.68" resultid="18623" heatid="19915" lane="4" entrytime="00:02:41.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="359" swimtime="00:01:10.07" resultid="18624" heatid="19978" lane="4" entrytime="00:01:10.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-07-04" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4823058" athleteid="18594">
              <RESULTS>
                <RESULT eventid="3551" points="352" swimtime="00:00:34.04" resultid="18595" heatid="19850" lane="6" entrytime="00:00:32.25" />
                <RESULT eventid="3649" points="426" reactiontime="+86" swimtime="00:02:15.55" resultid="18596" heatid="19896" lane="2" entrytime="00:02:12.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="427" swimtime="00:00:27.75" resultid="18597" heatid="19955" lane="6" entrytime="00:00:27.58" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-10-09" firstname="Julia3" gender="M" lastname="Janke-Frosch3" nation="ITA" swrid="4708009" athleteid="18598">
              <RESULTS>
                <RESULT eventid="3628" points="386" swimtime="00:01:20.43" resultid="18599" heatid="19870" lane="5" entrytime="00:01:19.58" />
                <RESULT eventid="3594" points="439" swimtime="00:00:27.50" resultid="18600" heatid="19954" lane="7" entrytime="00:00:28.01" />
                <RESULT eventid="3562" points="490" reactiontime="+82" swimtime="00:01:03.18" resultid="18601" heatid="19981" lane="8" entrytime="00:01:03.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-02-23" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4900633" athleteid="18561">
              <RESULTS>
                <RESULT eventid="3639" points="494" reactiontime="+70" swimtime="00:02:39.51" resultid="18562" heatid="19822" lane="8" entrytime="00:02:34.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="518" swimtime="00:01:20.21" resultid="18563" heatid="19862" lane="3" entrytime="00:01:19.90" />
                <RESULT eventid="3538" points="502" reactiontime="+66" swimtime="00:02:56.25" resultid="18564" heatid="19910" lane="6" entrytime="00:02:48.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-11-05" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4311786" athleteid="18516">
              <RESULTS>
                <RESULT eventid="3621" points="443" swimtime="00:01:24.54" resultid="18517" heatid="19861" lane="3" entrytime="00:01:22.89" />
                <RESULT eventid="3590" points="418" swimtime="00:00:31.73" resultid="18518" heatid="19929" lane="4" entrytime="00:00:31.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-02-04" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4911966" athleteid="18494">
              <RESULTS>
                <RESULT eventid="3621" points="237" swimtime="00:01:44.13" resultid="18495" heatid="19854" lane="4" entrytime="00:01:45.50" />
                <RESULT eventid="3570" points="268" swimtime="00:02:55.02" resultid="18496" heatid="19876" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-24" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4101995" athleteid="18532">
              <RESULTS>
                <RESULT eventid="3639" points="648" reactiontime="+42" swimtime="00:02:25.71" resultid="18533" heatid="19822" lane="4" entrytime="00:02:18.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="637" swimtime="00:02:11.28" resultid="18534" heatid="19888" lane="4" entrytime="00:02:04.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="637" reactiontime="+72" swimtime="00:01:05.12" resultid="18535" heatid="19975" lane="4" entrytime="00:00:59.99" />
                <RESULT eventid="3590" points="615" swimtime="00:00:27.90" resultid="19715" heatid="19936" lane="4" entrytime="00:00:26.30" />
                <RESULT eventid="15987" points="663" swimtime="00:00:27.21" resultid="20187" heatid="20132" lane="7" late="yes" />
                <RESULT eventid="15984" points="643" swimtime="00:00:27.48" resultid="20188" heatid="20130" lane="7" late="yes" />
                <RESULT eventid="15981" points="638" swimtime="00:00:27.56" resultid="20189" heatid="20128" lane="7" late="yes" />
                <RESULT eventid="15978" points="590" swimtime="00:00:28.29" resultid="20190" heatid="20126" lane="7" late="yes" />
                <RESULT eventid="15975" points="526" swimtime="00:00:29.38" resultid="20191" heatid="20124" lane="7" late="yes" />
                <RESULT eventid="15972" points="546" swimtime="00:00:29.03" resultid="20192" heatid="20122" lane="7" late="yes" />
                <RESULT eventid="15921" points="591" swimtime="00:00:28.27" resultid="20193" heatid="20120" lane="7" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-08-18" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4823063" athleteid="18508">
              <RESULTS>
                <RESULT eventid="3621" points="311" swimtime="00:01:35.12" resultid="18509" heatid="19856" lane="2" entrytime="00:01:40.05" />
                <RESULT eventid="3570" points="324" swimtime="00:02:44.47" resultid="18510" heatid="19879" lane="2" entrytime="00:02:51.12">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="329" swimtime="00:00:34.36" resultid="18511" heatid="19926" lane="6" entrytime="00:00:34.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-09-15" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4426768" athleteid="18569">
              <RESULTS>
                <RESULT eventid="3639" points="540" reactiontime="+80" swimtime="00:02:34.88" resultid="18570" heatid="19821" lane="6" entrytime="00:02:35.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="541" swimtime="00:00:29.11" resultid="18571" heatid="19936" lane="2" entrytime="00:00:28.80" />
                <RESULT eventid="3555" points="552" reactiontime="+78" swimtime="00:01:08.33" resultid="18572" heatid="19975" lane="6" entrytime="00:01:07.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-12-15" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4708010" athleteid="18649">
              <RESULTS>
                <RESULT eventid="3628" points="342" reactiontime="+70" swimtime="00:01:23.71" resultid="18650" heatid="19870" lane="6" entrytime="00:01:19.88" />
                <RESULT eventid="3594" points="369" swimtime="00:00:29.13" resultid="18651" heatid="19954" lane="3" entrytime="00:00:27.98" />
                <RESULT eventid="3562" points="389" reactiontime="+70" swimtime="00:01:08.21" resultid="18652" heatid="19980" lane="7" entrytime="00:01:06.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-06-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4823056" athleteid="18553">
              <RESULTS>
                <RESULT eventid="3621" points="393" reactiontime="+68" swimtime="00:01:27.95" resultid="18554" heatid="19861" lane="7" entrytime="00:01:23.90" />
                <RESULT eventid="3538" points="414" swimtime="00:03:07.94" resultid="18555" heatid="19908" lane="4" entrytime="00:03:00.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="382" swimtime="00:00:32.69" resultid="18556" heatid="19928" lane="4" entrytime="00:00:32.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-02-03" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4707986" athleteid="18501">
              <RESULTS>
                <RESULT eventid="3547" points="469" swimtime="00:00:34.82" resultid="18502" heatid="19843" lane="3" entrytime="00:00:33.90" />
                <RESULT eventid="3590" points="489" swimtime="00:00:30.10" resultid="18503" heatid="19934" lane="2" entrytime="00:00:29.98" />
                <RESULT eventid="3505" points="440" swimtime="00:02:44.04" resultid="18504" heatid="19993" lane="2" entrytime="00:02:30.12">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-10-22" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4823054" athleteid="18653">
              <RESULTS>
                <RESULT eventid="3628" points="207" reactiontime="+73" swimtime="00:01:39.01" resultid="18654" heatid="19867" lane="6" entrytime="00:01:30.12" />
                <RESULT eventid="3649" points="320" reactiontime="+49" swimtime="00:02:29.12" resultid="18655" heatid="19893" lane="3" entrytime="00:02:30.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-10" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4583010" athleteid="18645">
              <RESULTS>
                <RESULT eventid="3628" points="480" swimtime="00:01:14.79" resultid="18646" heatid="19871" lane="5" entrytime="00:01:14.56" />
                <RESULT eventid="3649" points="503" swimtime="00:02:08.23" resultid="18647" heatid="19898" lane="5" entrytime="00:02:03.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="470" reactiontime="+67" swimtime="00:02:43.65" resultid="18648" heatid="19916" lane="2" entrytime="00:02:32.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="423" swimtime="00:00:27.84" resultid="18658" heatid="19959" lane="1" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-02-18" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4800467" athleteid="18602">
              <RESULTS>
                <RESULT eventid="9711" points="669" reactiontime="+51" swimtime="00:02:10.33" resultid="18603" heatid="19832" lane="4" entrytime="00:02:03.36">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="620" swimtime="00:00:24.51" resultid="18604" heatid="19957" lane="4" entrytime="00:00:23.75" />
                <RESULT eventid="3562" points="645" reactiontime="+75" swimtime="00:00:57.64" resultid="18605" heatid="19982" lane="5" entrytime="00:00:57.88" />
                <RESULT eventid="15987" points="583" swimtime="00:00:25.03" resultid="20230" heatid="20133" lane="6" late="yes" />
                <RESULT eventid="15984" points="567" swimtime="00:00:25.25" resultid="20231" heatid="20131" lane="6" late="yes" />
                <RESULT eventid="15981" points="587" swimtime="00:00:24.96" resultid="20232" heatid="20129" lane="6" late="yes" />
                <RESULT eventid="15978" points="587" swimtime="00:00:24.97" resultid="20233" heatid="20127" lane="6" late="yes" />
                <RESULT eventid="15975" points="555" swimtime="00:00:25.44" resultid="20234" heatid="20125" lane="6" late="yes" />
                <RESULT eventid="15972" points="557" swimtime="00:00:25.41" resultid="20235" heatid="20123" lane="6" late="yes" />
                <RESULT eventid="15921" points="587" swimtime="00:00:24.96" resultid="20236" heatid="20121" lane="6" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-10-27" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4911971" athleteid="18606">
              <RESULTS>
                <RESULT eventid="3649" points="323" swimtime="00:02:28.57" resultid="18607" heatid="19891" lane="5" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="275" swimtime="00:00:32.12" resultid="18608" heatid="19950" lane="8" entrytime="00:00:34.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-04-09" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4823066" athleteid="18528">
              <RESULTS>
                <RESULT eventid="3639" points="428" swimtime="00:02:47.30" resultid="18529" heatid="19818" lane="3" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="427" swimtime="00:00:35.91" resultid="18530" heatid="19842" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="3505" points="443" swimtime="00:02:43.71" resultid="18531" heatid="19991" lane="8" entrytime="00:02:40.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-05-19" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4708011" athleteid="18577">
              <RESULTS>
                <RESULT eventid="3621" points="453" reactiontime="+74" swimtime="00:01:23.89" resultid="18578" heatid="19861" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="3570" points="479" reactiontime="+78" swimtime="00:02:24.37" resultid="18579" heatid="19885" lane="6" entrytime="00:02:23.65">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="404" swimtime="00:03:09.43" resultid="18580" heatid="19909" lane="3" entrytime="00:02:53.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="426" swimtime="00:00:31.52" resultid="18581" heatid="19931" lane="5" entrytime="00:00:30.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-12-07" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4707988" athleteid="18625">
              <RESULTS>
                <RESULT eventid="9711" points="522" swimtime="00:02:21.58" resultid="18626" heatid="19831" lane="4" entrytime="00:02:21.12">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="478" swimtime="00:00:30.73" resultid="18627" heatid="19851" lane="5" entrytime="00:00:30.08" />
                <RESULT eventid="3512" points="525" swimtime="00:02:18.67" resultid="18628" heatid="20001" lane="5" entrytime="00:02:13.32">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-04-02" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4823061" athleteid="18633">
              <RESULTS>
                <RESULT eventid="9711" points="398" swimtime="00:02:34.88" resultid="18634" heatid="19830" lane="3" entrytime="00:02:29.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="415" swimtime="00:00:32.21" resultid="18635" heatid="19850" lane="7" entrytime="00:00:32.56" />
                <RESULT eventid="3512" points="435" swimtime="00:02:27.60" resultid="18636" heatid="20001" lane="7" entrytime="00:02:20.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-02-04" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5150855" athleteid="18512">
              <RESULTS>
                <RESULT eventid="3547" points="448" swimtime="00:00:35.34" resultid="18513" heatid="19842" lane="1" entrytime="00:00:36.01" />
                <RESULT eventid="3590" points="421" swimtime="00:00:31.65" resultid="18514" heatid="19929" lane="1" entrytime="00:00:32.22" />
                <RESULT eventid="3505" points="363" swimtime="00:02:54.91" resultid="18515" heatid="19989" lane="4" entrytime="00:02:45.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-09-27" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4708025" athleteid="18586">
              <RESULTS>
                <RESULT eventid="3639" points="518" swimtime="00:02:37.02" resultid="18587" heatid="19822" lane="2" entrytime="00:02:30.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="544" reactiontime="+70" swimtime="00:02:18.39" resultid="18588" heatid="19888" lane="1" entrytime="00:02:13.89">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="470" swimtime="00:02:40.49" resultid="18589" heatid="19992" lane="6" entrytime="00:02:33.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-11-26" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4708001" athleteid="18519">
              <RESULTS>
                <RESULT eventid="3547" points="426" swimtime="00:00:35.95" resultid="18520" heatid="19843" lane="8" entrytime="00:00:34.80" />
                <RESULT eventid="3570" points="427" reactiontime="+50" swimtime="00:02:30.01" resultid="18521" heatid="19883" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="394" swimtime="00:02:50.16" resultid="18522" heatid="19992" lane="1" entrytime="00:02:36.65">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-04-03" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5089281" athleteid="18582">
              <RESULTS>
                <RESULT eventid="3547" points="273" swimtime="00:00:41.69" resultid="18583" heatid="19839" lane="4" entrytime="00:00:40.10" />
                <RESULT eventid="3590" points="250" swimtime="00:00:37.62" resultid="18584" heatid="19925" lane="7" entrytime="00:00:35.40" />
                <RESULT eventid="3505" points="269" swimtime="00:03:13.24" resultid="18585" heatid="19985" lane="3" entrytime="00:03:09.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-08-29" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4929228" athleteid="18549">
              <RESULTS>
                <RESULT eventid="3639" points="495" reactiontime="+93" swimtime="00:02:39.45" resultid="18550" heatid="19819" lane="7" entrytime="00:02:42.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="497" reactiontime="+77" swimtime="00:01:21.34" resultid="18551" heatid="19862" lane="6" entrytime="00:01:20.50" />
                <RESULT eventid="3538" points="480" swimtime="00:02:58.90" resultid="18552" heatid="19909" lane="5" entrytime="00:02:52.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="12820" points="474" swimtime="00:04:25.70" resultid="18660" heatid="20141" lane="7" entrytime="00:04:20.16">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="200" swimtime="00:02:22.41" />
                    <SPLIT distance="300" swimtime="00:03:26.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18625" number="1" />
                    <RELAYPOSITION athleteid="18621" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="18598" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="18613" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="3574" points="490" swimtime="00:04:54.44" resultid="18659" heatid="20139" lane="3" entrytime="00:04:44.16">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="200" swimtime="00:02:39.69" />
                    <SPLIT distance="300" swimtime="00:03:47.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18512" number="1" />
                    <RELAYPOSITION athleteid="18549" number="2" reactiontime="+6" />
                    <RELAYPOSITION athleteid="18569" number="3" reactiontime="+12" />
                    <RELAYPOSITION athleteid="18565" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MIH" nation="AUT" region="TLSV" clubid="16577" swrid="89762" name="Breedy Badger" shortname="MIH Zillertal">
          <CONTACT city="Bruck am Ziller" email="swim@make-it-happen.at" internet="www.make-it-happen.at" name="Breedy Badger" phone="06769734383" state="TI" street="Dorf 42d" zip="6260" />
          <ATHLETES>
            <ATHLETE birthdate="2005-05-04" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43378" swrid="4953384" athleteid="16587">
              <RESULTS>
                <RESULT eventid="3639" points="326" swimtime="00:03:03.14" resultid="16588" heatid="19815" lane="6" entrytime="00:02:57.32">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="319" swimtime="00:01:34.24" resultid="16589" heatid="19858" lane="7" entrytime="00:01:34.08" />
                <RESULT eventid="3570" points="352" swimtime="00:02:40.00" resultid="16590" heatid="19881" lane="6" entrytime="00:02:38.12">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="320" swimtime="00:01:21.93" resultid="16591" heatid="19971" lane="7" entrytime="00:01:21.26" />
                <RESULT eventid="3505" points="345" swimtime="00:02:57.82" resultid="16592" heatid="19989" lane="1" entrytime="00:02:50.22">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="368" swimtime="00:01:21.09" resultid="16593" heatid="20009" lane="2" entrytime="00:01:18.45" />
                <RESULT eventid="3658" points="321" swimtime="00:05:49.24" resultid="16594" heatid="20045" lane="1" entrytime="00:05:34.21">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.07" />
                    <SPLIT distance="200" swimtime="00:02:52.12" />
                    <SPLIT distance="300" swimtime="00:04:24.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="382" swimtime="00:01:11.74" resultid="16595" heatid="20091" lane="4" entrytime="00:01:11.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-14" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="42402" swrid="5029804" athleteid="16596">
              <RESULTS>
                <RESULT eventid="9711" points="240" swimtime="00:03:03.39" resultid="16597" heatid="19827" lane="2" entrytime="00:02:52.26">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="186" swimtime="00:01:42.50" resultid="16598" heatid="19865" lane="5" entrytime="00:01:36.24" />
                <RESULT eventid="3649" points="248" reactiontime="+51" swimtime="00:02:42.19" resultid="16599" heatid="19893" lane="7" entrytime="00:02:34.60">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="163" reactiontime="+55" swimtime="00:01:31.12" resultid="16600" heatid="19977" lane="6" entrytime="00:01:21.79" />
                <RESULT eventid="3512" points="245" swimtime="00:02:58.86" resultid="16601" heatid="19998" lane="7" entrytime="00:02:47.31">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="219" swimtime="00:01:26.14" resultid="16602" heatid="20017" lane="6" entrytime="00:01:19.38" />
                <RESULT eventid="3578" points="273" reactiontime="+48" swimtime="00:05:39.04" resultid="16603" heatid="20055" lane="8" entrytime="00:05:29.83">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="200" swimtime="00:02:47.80" />
                    <SPLIT distance="300" swimtime="00:04:14.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="249" reactiontime="+57" swimtime="00:01:14.56" resultid="16604" heatid="20105" lane="1" entrytime="00:01:11.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-10-27" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42622" swrid="5055504" athleteid="16578">
              <RESULTS>
                <RESULT eventid="3639" points="380" reactiontime="+76" swimtime="00:02:54.14" resultid="16579" heatid="19818" lane="7" entrytime="00:02:46.79">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="300" reactiontime="+71" swimtime="00:01:36.27" resultid="16580" heatid="19858" lane="1" entrytime="00:01:34.27" />
                <RESULT eventid="3570" points="419" swimtime="00:02:30.95" resultid="16581" heatid="19883" lane="8" entrytime="00:02:30.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="391" swimtime="00:01:16.66" resultid="16582" heatid="19971" lane="4" entrytime="00:01:19.38" />
                <RESULT eventid="3505" points="392" swimtime="00:02:50.47" resultid="16583" heatid="19990" lane="5" entrytime="00:02:42.05">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="375" swimtime="00:01:20.57" resultid="16584" heatid="20009" lane="6" entrytime="00:01:18.06" />
                <RESULT eventid="3658" points="417" swimtime="00:05:19.90" resultid="16585" heatid="20046" lane="3" entrytime="00:05:12.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.55" />
                    <SPLIT distance="200" swimtime="00:02:37.84" />
                    <SPLIT distance="300" swimtime="00:04:00.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="413" reactiontime="+82" swimtime="00:01:09.89" resultid="16586" heatid="20093" lane="6" entrytime="00:01:09.15" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RARINANT" nation="ITA" clubid="17497" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5006758" athleteid="17819">
              <RESULTS>
                <RESULT eventid="3621" points="316" reactiontime="+67" swimtime="00:01:34.58" resultid="17820" heatid="19857" lane="7" entrytime="00:01:36.66" />
                <RESULT eventid="3538" points="335" swimtime="00:03:21.73" resultid="17821" heatid="19905" lane="5" entrytime="00:03:34.51">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="277" swimtime="00:01:29.11" resultid="17822" heatid="20003" lane="4" entrytime="00:01:33.68" />
                <RESULT eventid="3523" points="323" reactiontime="+76" swimtime="00:01:15.86" resultid="17823" heatid="20087" lane="6" entrytime="00:01:20.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4938672" athleteid="17841">
              <RESULTS>
                <RESULT eventid="3621" points="354" swimtime="00:01:31.09" resultid="17842" heatid="19857" lane="5" entrytime="00:01:35.00" />
                <RESULT eventid="3505" points="319" swimtime="00:03:02.60" resultid="17843" heatid="19986" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="345" reactiontime="+64" swimtime="00:05:40.92" resultid="17844" heatid="20045" lane="8" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.29" />
                    <SPLIT distance="200" swimtime="00:02:45.32" />
                    <SPLIT distance="300" swimtime="00:04:13.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4585060" athleteid="17706">
              <RESULTS>
                <RESULT eventid="3551" points="505" swimtime="00:00:30.17" resultid="17707" heatid="19851" lane="4" entrytime="00:00:29.90" />
                <RESULT eventid="3512" points="531" swimtime="00:02:18.20" resultid="17708" heatid="20001" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="527" swimtime="00:01:04.30" resultid="17709" heatid="20022" lane="1" entrytime="00:01:03.50" />
                <RESULT eventid="3613" points="458" swimtime="00:00:29.08" resultid="17710" heatid="20037" lane="5" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4500996" athleteid="17696">
              <RESULTS>
                <RESULT eventid="3649" points="496" reactiontime="+66" swimtime="00:02:08.78" resultid="17697" heatid="19898" lane="2" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="483" reactiontime="+66" swimtime="00:01:03.47" resultid="17698" heatid="19981" lane="2" entrytime="00:01:02.80" />
                <RESULT eventid="3605" points="427" swimtime="00:01:08.94" resultid="17699" heatid="20020" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="3588" points="469" reactiontime="+68" swimtime="00:02:23.43" resultid="17700" heatid="20067" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4907158" athleteid="17507">
              <RESULTS>
                <RESULT eventid="3639" points="350" swimtime="00:02:58.89" resultid="17508" heatid="19813" lane="3" entrytime="00:03:04.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="422" swimtime="00:00:31.63" resultid="17509" heatid="19931" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="3523" points="461" swimtime="00:01:07.39" resultid="17510" heatid="20094" lane="5" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4504630" athleteid="17768">
              <RESULTS>
                <RESULT eventid="3547" points="529" swimtime="00:00:33.45" resultid="17769" heatid="19843" lane="5" entrytime="00:00:33.54" />
                <RESULT eventid="3555" points="555" reactiontime="+83" swimtime="00:01:08.21" resultid="17770" heatid="19974" lane="4" entrytime="00:01:08.61" />
                <RESULT eventid="3617" points="562" swimtime="00:00:30.37" resultid="17771" heatid="20031" lane="1" entrytime="00:00:30.42" />
                <RESULT eventid="3523" points="484" reactiontime="+79" swimtime="00:01:06.29" resultid="17772" heatid="20096" lane="4" entrytime="00:01:05.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4843909" athleteid="17758">
              <RESULTS>
                <RESULT eventid="9711" points="435" swimtime="00:02:30.38" resultid="17759" heatid="19830" lane="5" entrytime="00:02:29.42">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="436" reactiontime="+67" swimtime="00:02:14.48" resultid="17760" heatid="19895" lane="2" entrytime="00:02:16.88">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="342" swimtime="00:01:14.27" resultid="17761" heatid="20018" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1081" points="431" swimtime="00:05:22.75" resultid="17762" heatid="20118" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="200" swimtime="00:02:40.57" />
                    <SPLIT distance="300" swimtime="00:04:09.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4809373" athleteid="17631">
              <RESULTS>
                <RESULT eventid="3649" points="371" reactiontime="+52" swimtime="00:02:21.85" resultid="17632" heatid="19896" lane="8" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="357" swimtime="00:00:29.45" resultid="17633" heatid="19952" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="3613" points="334" swimtime="00:00:32.30" resultid="17634" heatid="20036" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="3530" points="361" reactiontime="+63" swimtime="00:01:05.86" resultid="17635" heatid="20108" lane="2" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4717997" athleteid="17558">
              <RESULTS>
                <RESULT eventid="3570" points="557" reactiontime="+76" swimtime="00:02:17.28" resultid="17559" heatid="19888" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="618" swimtime="00:00:27.85" resultid="17560" heatid="19935" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="3617" points="548" swimtime="00:00:30.62" resultid="17561" heatid="20031" lane="7" entrytime="00:00:30.30" />
                <RESULT eventid="3523" points="594" reactiontime="+64" swimtime="00:01:01.93" resultid="17562" heatid="20099" lane="4" entrytime="00:00:59.98" />
                <RESULT eventid="15921" points="620" swimtime="00:00:27.82" resultid="20180" heatid="20120" lane="2" late="yes" />
                <RESULT eventid="15972" points="526" swimtime="00:00:29.39" resultid="20181" heatid="20122" lane="2" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4695537" athleteid="17726">
              <RESULTS>
                <RESULT eventid="3628" points="499" reactiontime="+87" swimtime="00:01:13.83" resultid="17727" heatid="19871" lane="6" entrytime="00:01:15.99" />
                <RESULT eventid="3545" points="491" reactiontime="+78" swimtime="00:02:41.34" resultid="17728" heatid="19916" lane="8" entrytime="00:02:40.76">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="452" swimtime="00:01:07.66" resultid="17729" heatid="20020" lane="4" entrytime="00:01:08.34" />
                <RESULT eventid="1081" points="515" reactiontime="+69" swimtime="00:05:04.19" resultid="17730" heatid="20119" lane="6" entrytime="00:04:56.81">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.77" />
                    <SPLIT distance="200" swimtime="00:02:26.57" />
                    <SPLIT distance="300" swimtime="00:03:53.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4929528" athleteid="17586">
              <RESULTS>
                <RESULT eventid="3628" points="200" reactiontime="+71" swimtime="00:01:40.07" resultid="17587" heatid="19866" lane="7" entrytime="00:01:34.55" />
                <RESULT eventid="3512" points="298" swimtime="00:02:47.50" resultid="17588" heatid="19998" lane="1" entrytime="00:02:47.71">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="304" reactiontime="+63" swimtime="00:05:27.25" resultid="17589" heatid="20055" lane="1" entrytime="00:05:28.48">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.24" />
                    <SPLIT distance="200" swimtime="00:02:42.15" />
                    <SPLIT distance="300" swimtime="00:04:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="265" reactiontime="+61" swimtime="00:06:19.54" resultid="17590" heatid="20117" lane="1" entrytime="00:06:10.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                    <SPLIT distance="200" swimtime="00:03:03.71" />
                    <SPLIT distance="300" swimtime="00:04:58.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" athleteid="17833">
              <RESULTS>
                <RESULT eventid="3639" points="384" reactiontime="+64" swimtime="00:02:53.52" resultid="17834" heatid="19816" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="344" swimtime="00:02:57.99" resultid="17835" heatid="19987" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="395" swimtime="00:01:10.95" resultid="17836" heatid="20093" lane="8" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5006757" athleteid="17798">
              <RESULTS>
                <RESULT eventid="3621" points="465" reactiontime="+55" swimtime="00:01:23.18" resultid="17799" heatid="19862" lane="8" entrytime="00:01:22.00" />
                <RESULT eventid="3590" points="372" swimtime="00:00:32.98" resultid="17800" heatid="19925" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="3586" points="340" swimtime="00:02:54.39" resultid="17801" heatid="20063" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5039265" athleteid="17802">
              <RESULTS>
                <RESULT eventid="3555" status="DNS" swimtime="00:00:00.00" resultid="17803" heatid="19970" lane="5" entrytime="00:01:25.00" />
                <RESULT eventid="3598" points="279" swimtime="00:01:28.94" resultid="17804" heatid="20006" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="3523" points="365" reactiontime="+63" swimtime="00:01:12.80" resultid="17805" heatid="20094" lane="4" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="5176663" athleteid="17498">
              <RESULTS>
                <RESULT eventid="3649" points="207" swimtime="00:02:52.32" resultid="17499" heatid="19890" lane="5" entrytime="00:02:50.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="219" swimtime="00:03:05.53" resultid="17500" heatid="19997" lane="2" entrytime="00:02:57.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="227" swimtime="00:06:00.41" resultid="17501" heatid="20053" lane="4" entrytime="00:05:43.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.27" />
                    <SPLIT distance="200" swimtime="00:02:57.79" />
                    <SPLIT distance="300" swimtime="00:04:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="207" reactiontime="+74" swimtime="00:01:19.22" resultid="17502" heatid="20101" lane="7" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4500981" athleteid="17850">
              <RESULTS>
                <RESULT eventid="3570" points="480" reactiontime="+70" swimtime="00:02:24.23" resultid="17851" heatid="19886" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment=" - Hat den Wettkampf nicht in der gleichen Bahn beendet (Zeit: 17:18)" eventid="3505" status="DSQ" swimtime="00:02:44.89" resultid="17852" heatid="19992" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3617" points="367" swimtime="00:00:35.01" resultid="17853" heatid="20028" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="3523" points="456" reactiontime="+87" swimtime="00:01:07.62" resultid="17854" heatid="20097" lane="5" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4843914" athleteid="17744">
              <RESULTS>
                <RESULT eventid="3562" points="321" reactiontime="+79" swimtime="00:01:12.69" resultid="17745" heatid="19978" lane="8" entrytime="00:01:18.54" />
                <RESULT eventid="3578" points="464" reactiontime="+74" swimtime="00:04:44.15" resultid="17746" heatid="20057" lane="7" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.80" />
                    <SPLIT distance="200" swimtime="00:02:19.09" />
                    <SPLIT distance="300" swimtime="00:03:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3588" points="307" reactiontime="+85" swimtime="00:02:45.14" resultid="17747" heatid="20066" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="403" reactiontime="+64" swimtime="00:01:03.46" resultid="17748" heatid="20107" lane="3" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4641186" athleteid="17606">
              <RESULTS>
                <RESULT eventid="9711" points="421" reactiontime="+74" swimtime="00:02:32.03" resultid="17607" heatid="19830" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="372" swimtime="00:00:29.05" resultid="17608" heatid="19954" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="3578" points="427" reactiontime="+67" swimtime="00:04:52.23" resultid="17609" heatid="20057" lane="1" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.08" />
                    <SPLIT distance="200" swimtime="00:02:20.66" />
                    <SPLIT distance="300" swimtime="00:03:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3588" points="418" reactiontime="+70" swimtime="00:02:29.09" resultid="17610" heatid="20067" lane="6" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4929529" athleteid="17829">
              <RESULTS>
                <RESULT eventid="3555" points="350" swimtime="00:01:19.48" resultid="17830" heatid="19971" lane="3" entrytime="00:01:20.00" />
                <RESULT eventid="3658" points="428" swimtime="00:05:17.29" resultid="17831" heatid="20046" lane="2" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.28" />
                    <SPLIT distance="200" swimtime="00:02:34.86" />
                    <SPLIT distance="300" swimtime="00:03:56.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3636" points="440" reactiontime="+62" swimtime="00:05:54.04" resultid="17832" heatid="20114" lane="6" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                    <SPLIT distance="200" swimtime="00:02:55.53" />
                    <SPLIT distance="300" swimtime="00:04:32.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4907157" athleteid="17591">
              <RESULTS>
                <RESULT eventid="3570" points="449" reactiontime="+91" swimtime="00:02:27.48" resultid="17592" heatid="19884" lane="6" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="408" swimtime="00:00:31.97" resultid="17593" heatid="19930" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="3658" points="465" swimtime="00:05:08.48" resultid="17594" heatid="20046" lane="5" entrytime="00:05:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.10" />
                    <SPLIT distance="200" swimtime="00:02:32.21" />
                    <SPLIT distance="300" swimtime="00:03:51.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="427" reactiontime="+81" swimtime="00:01:09.10" resultid="17595" heatid="20093" lane="7" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4695607" athleteid="17731">
              <RESULTS>
                <RESULT eventid="3594" points="483" swimtime="00:00:26.64" resultid="17732" heatid="19956" lane="2" entrytime="00:00:27.18" />
                <RESULT eventid="3605" points="476" swimtime="00:01:06.51" resultid="17733" heatid="20021" lane="5" entrytime="00:01:04.99" />
                <RESULT eventid="3578" points="527" reactiontime="+70" swimtime="00:04:32.31" resultid="17734" heatid="20057" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.71" />
                    <SPLIT distance="200" swimtime="00:02:13.40" />
                    <SPLIT distance="300" swimtime="00:03:24.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="546" reactiontime="+70" swimtime="00:00:57.37" resultid="17735" heatid="20110" lane="8" entrytime="00:00:59.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4586112" athleteid="17691">
              <RESULTS>
                <RESULT eventid="3628" points="693" swimtime="00:01:06.19" resultid="17692" heatid="19872" lane="5" entrytime="00:01:05.50" />
                <RESULT eventid="3545" points="577" reactiontime="+52" swimtime="00:02:32.91" resultid="17693" heatid="19916" lane="3" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3613" points="479" swimtime="00:00:28.65" resultid="17694" heatid="20038" lane="2" entrytime="00:00:28.80" />
                <RESULT eventid="3519" points="627" swimtime="00:00:31.15" resultid="17695" heatid="20084" lane="4" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4695535" athleteid="17721">
              <RESULTS>
                <RESULT comment=" - Delphinkick nach jedem Brustbeinschlag (Zeit: 12:46)" eventid="3628" reactiontime="+58" status="DSQ" swimtime="00:01:15.03" resultid="17722" heatid="19870" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="3562" points="505" reactiontime="+62" swimtime="00:01:02.56" resultid="17723" heatid="19981" lane="5" entrytime="00:01:02.00" />
                <RESULT eventid="3605" points="394" swimtime="00:01:10.79" resultid="17724" heatid="20018" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="3588" points="476" reactiontime="+67" swimtime="00:02:22.79" resultid="17725" heatid="20067" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="5006998" athleteid="17666">
              <RESULTS>
                <RESULT eventid="3628" points="214" reactiontime="+78" swimtime="00:01:37.91" resultid="17667" heatid="19865" lane="6" entrytime="00:01:37.16" />
                <RESULT eventid="3562" points="267" swimtime="00:01:17.28" resultid="17668" heatid="19977" lane="2" entrytime="00:01:22.00" />
                <RESULT eventid="3605" points="296" swimtime="00:01:17.92" resultid="17669" heatid="20017" lane="4" entrytime="00:01:18.11" />
                <RESULT eventid="1081" points="281" swimtime="00:06:11.88" resultid="17670" heatid="20117" lane="8" entrytime="00:06:13.03">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.62" />
                    <SPLIT distance="200" swimtime="00:02:55.89" />
                    <SPLIT distance="300" swimtime="00:04:47.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" athleteid="17763">
              <RESULTS>
                <RESULT eventid="9711" points="531" reactiontime="+60" swimtime="00:02:20.70" resultid="17764" heatid="19832" lane="7" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="547" reactiontime="+49" swimtime="00:01:00.90" resultid="17765" heatid="19982" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="3613" points="567" swimtime="00:00:27.09" resultid="17766" heatid="20039" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="3530" points="566" reactiontime="+62" swimtime="00:00:56.70" resultid="17767" heatid="20111" lane="2" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4907159" athleteid="17511">
              <RESULTS>
                <RESULT eventid="3547" points="227" swimtime="00:00:44.33" resultid="17512" heatid="19838" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="3590" points="313" swimtime="00:00:34.95" resultid="17513" heatid="19924" lane="4" entrytime="00:00:35.80" />
                <RESULT eventid="3523" points="283" reactiontime="+69" swimtime="00:01:19.22" resultid="17514" heatid="20086" lane="4" entrytime="00:01:24.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5124159" athleteid="17661">
              <RESULTS>
                <RESULT eventid="3621" points="206" reactiontime="+57" swimtime="00:01:49.11" resultid="17662" heatid="19854" lane="7" entrytime="00:01:48.38" />
                <RESULT eventid="3505" points="322" swimtime="00:03:01.95" resultid="17663" heatid="19988" lane="5" entrytime="00:02:52.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="324" swimtime="00:01:24.54" resultid="17664" heatid="20008" lane="6" entrytime="00:01:20.70" />
                <RESULT eventid="3658" points="317" reactiontime="+55" swimtime="00:05:50.62" resultid="17665" heatid="20041" lane="6" entrytime="00:06:18.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.79" />
                    <SPLIT distance="200" swimtime="00:02:51.93" />
                    <SPLIT distance="300" swimtime="00:04:22.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5001363" athleteid="17515">
              <RESULTS>
                <RESULT eventid="3639" points="317" reactiontime="+75" swimtime="00:03:04.84" resultid="17516" heatid="19814" lane="1" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="316" swimtime="00:03:25.71" resultid="17517" heatid="19906" lane="4" entrytime="00:03:25.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="324" swimtime="00:00:43.38" resultid="17518" heatid="20071" lane="4" entrytime="00:00:44.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4750725" athleteid="17616">
              <RESULTS>
                <RESULT eventid="3649" points="391" swimtime="00:02:19.48" resultid="17617" heatid="19896" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="399" swimtime="00:00:28.40" resultid="17618" heatid="19953" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="3613" points="355" swimtime="00:00:31.67" resultid="17619" heatid="20036" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="3588" points="334" reactiontime="+82" swimtime="00:02:40.71" resultid="17620" heatid="20067" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4809440" athleteid="17601">
              <RESULTS>
                <RESULT eventid="3628" points="429" reactiontime="+66" swimtime="00:01:17.66" resultid="17602" heatid="19869" lane="4" entrytime="00:01:20.00" />
                <RESULT eventid="3545" points="397" reactiontime="+74" swimtime="00:02:53.16" resultid="17603" heatid="19915" lane="8" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3613" points="281" swimtime="00:00:34.24" resultid="17604" heatid="20035" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="3519" points="437" swimtime="00:00:35.14" resultid="17605" heatid="20082" lane="4" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4809382" athleteid="17621">
              <RESULTS>
                <RESULT eventid="3649" points="351" reactiontime="+68" swimtime="00:02:24.54" resultid="17622" heatid="19896" lane="7" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="386" reactiontime="+71" swimtime="00:01:08.38" resultid="17623" heatid="19980" lane="8" entrytime="00:01:07.00" />
                <RESULT eventid="3613" points="415" swimtime="00:00:30.07" resultid="17624" heatid="20036" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="3530" status="DNS" swimtime="00:00:00.00" resultid="17625" heatid="20108" lane="7" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4938680" athleteid="17837">
              <RESULTS>
                <RESULT eventid="3639" points="336" swimtime="00:03:01.40" resultid="17838" heatid="19814" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="339" swimtime="00:05:42.76" resultid="17839" heatid="20042" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="200" swimtime="00:02:48.64" />
                    <SPLIT distance="300" swimtime="00:04:17.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="343" reactiontime="+58" swimtime="00:01:14.33" resultid="17840" heatid="20090" lane="1" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4495015" athleteid="17543">
              <RESULTS>
                <RESULT eventid="3547" points="602" swimtime="00:00:32.04" resultid="17544" heatid="19844" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="3590" points="492" swimtime="00:00:30.05" resultid="17545" heatid="19935" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="3598" status="DNS" swimtime="00:00:00.00" resultid="17546" heatid="20012" lane="4" entrytime="00:01:09.50" />
                <RESULT eventid="3523" status="DNS" swimtime="00:00:00.00" resultid="17547" heatid="20098" lane="7" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4843901" athleteid="17754">
              <RESULTS>
                <RESULT eventid="3628" points="407" swimtime="00:01:19.03" resultid="17755" heatid="19869" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="3562" points="419" reactiontime="+47" swimtime="00:01:06.54" resultid="17756" heatid="19980" lane="1" entrytime="00:01:07.00" />
                <RESULT eventid="3530" points="374" reactiontime="+43" swimtime="00:01:05.10" resultid="17757" heatid="20107" lane="5" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4907162" athleteid="17519">
              <RESULTS>
                <RESULT eventid="3649" points="384" swimtime="00:02:20.28" resultid="17520" heatid="19894" lane="3" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="337" swimtime="00:01:11.58" resultid="17521" heatid="19979" lane="1" entrytime="00:01:09.00" />
                <RESULT eventid="1081" points="350" swimtime="00:05:45.77" resultid="17522" heatid="20117" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="200" swimtime="00:02:51.84" />
                    <SPLIT distance="300" swimtime="00:04:31.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4500971" athleteid="17845">
              <RESULTS>
                <RESULT eventid="3570" points="612" swimtime="00:02:13.02" resultid="17846" heatid="19888" lane="5" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="619" swimtime="00:00:27.84" resultid="17847" heatid="19936" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="3658" points="587" reactiontime="+71" swimtime="00:04:45.46" resultid="17848" heatid="20050" lane="2" entrytime="00:04:43.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="200" swimtime="00:02:16.97" />
                    <SPLIT distance="300" swimtime="00:03:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="434" swimtime="00:00:39.34" resultid="17849" heatid="20075" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="15978" points="557" swimtime="00:00:28.83" resultid="20176" heatid="20126" lane="6" late="yes" />
                <RESULT eventid="15975" points="532" swimtime="00:00:29.27" resultid="20177" heatid="20124" lane="6" late="yes" />
                <RESULT eventid="15972" points="549" swimtime="00:00:28.97" resultid="20178" heatid="20122" lane="6" late="yes" />
                <RESULT eventid="15921" points="593" swimtime="00:00:28.24" resultid="20179" heatid="20120" lane="6" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4809381" athleteid="17626">
              <RESULTS>
                <RESULT eventid="3649" points="498" reactiontime="+57" swimtime="00:02:08.66" resultid="17627" heatid="19898" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="482" swimtime="00:00:26.66" resultid="17628" heatid="19957" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="3605" points="431" swimtime="00:01:08.72" resultid="17629" heatid="20020" lane="7" entrytime="00:01:11.00" />
                <RESULT eventid="3530" points="506" reactiontime="+72" swimtime="00:00:58.85" resultid="17630" heatid="20111" lane="1" entrytime="00:00:56.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4907161" athleteid="17527">
              <RESULTS>
                <RESULT eventid="3649" points="375" reactiontime="+77" swimtime="00:02:21.34" resultid="17528" heatid="19894" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="364" swimtime="00:02:36.73" resultid="17529" heatid="19999" lane="3" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="369" reactiontime="+73" swimtime="00:01:05.35" resultid="17530" heatid="20107" lane="2" entrytime="00:01:06.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5039263" athleteid="17646">
              <RESULTS>
                <RESULT eventid="3570" points="309" swimtime="00:02:47.02" resultid="17647" heatid="19876" lane="3" entrytime="00:03:02.88">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="240" swimtime="00:03:20.76" resultid="17648" heatid="19986" lane="3" entrytime="00:03:04.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="296" reactiontime="+57" swimtime="00:05:58.52" resultid="17649" heatid="20042" lane="7" entrytime="00:06:08.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="200" swimtime="00:02:59.32" />
                    <SPLIT distance="300" swimtime="00:04:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="253" swimtime="00:01:22.28" resultid="17650" heatid="20089" lane="8" entrytime="00:01:16.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5006993" athleteid="17656">
              <RESULTS>
                <RESULT eventid="3570" points="301" swimtime="00:02:48.53" resultid="17657" heatid="19878" lane="5" entrytime="00:02:54.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="253" swimtime="00:01:28.59" resultid="17658" heatid="19968" lane="5" entrytime="00:01:35.94" />
                <RESULT eventid="3598" points="252" swimtime="00:01:31.92" resultid="17659" heatid="20004" lane="6" entrytime="00:01:32.00" />
                <RESULT eventid="3636" points="347" swimtime="00:06:23.18" resultid="17660" heatid="20114" lane="8" entrytime="00:06:18.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.12" />
                    <SPLIT distance="200" swimtime="00:03:08.52" />
                    <SPLIT distance="300" swimtime="00:04:55.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4585058" athleteid="17783">
              <RESULTS>
                <RESULT eventid="3570" points="422" reactiontime="+66" swimtime="00:02:30.55" resultid="17784" heatid="19884" lane="2" entrytime="00:02:26.24">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="366" swimtime="00:00:33.16" resultid="17785" heatid="19932" lane="8" entrytime="00:00:30.84" />
                <RESULT eventid="3598" points="321" swimtime="00:01:24.82" resultid="17786" heatid="20006" lane="1" entrytime="00:01:26.30" />
                <RESULT eventid="3586" points="353" swimtime="00:02:52.29" resultid="17787" heatid="20065" lane="8" entrytime="00:02:42.17">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4641072" athleteid="17701">
              <RESULTS>
                <RESULT eventid="3628" points="594" reactiontime="+83" swimtime="00:01:09.66" resultid="17702" heatid="19872" lane="2" entrytime="00:01:10.00" />
                <RESULT eventid="3545" points="611" reactiontime="+84" swimtime="00:02:29.98" resultid="17703" heatid="19916" lane="6" entrytime="00:02:30.95">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="615" reactiontime="+79" swimtime="00:04:18.71" resultid="17704" heatid="20058" lane="2" entrytime="00:04:21.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.57" />
                    <SPLIT distance="200" swimtime="00:02:08.06" />
                    <SPLIT distance="300" swimtime="00:03:15.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="588" reactiontime="+74" swimtime="00:04:50.92" resultid="17705" heatid="20119" lane="3" entrytime="00:04:52.51">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.16" />
                    <SPLIT distance="200" swimtime="00:02:27.60" />
                    <SPLIT distance="300" swimtime="00:03:45.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" athleteid="17711">
              <RESULTS>
                <RESULT eventid="9711" points="478" reactiontime="+61" swimtime="00:02:25.80" resultid="17712" heatid="19831" lane="7" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="459" swimtime="00:00:27.09" resultid="17713" heatid="19955" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="3562" points="488" reactiontime="+54" swimtime="00:01:03.24" resultid="17714" heatid="19980" lane="4" entrytime="00:01:03.50" />
                <RESULT eventid="3613" points="498" swimtime="00:00:28.28" resultid="17715" heatid="20038" lane="6" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4843906" athleteid="17824">
              <RESULTS>
                <RESULT eventid="3639" points="389" reactiontime="+78" swimtime="00:02:52.77" resultid="17825" heatid="19814" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="412" swimtime="00:02:47.70" resultid="17826" heatid="19990" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="464" reactiontime="+80" swimtime="00:05:08.69" resultid="17827" heatid="20047" lane="7" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="200" swimtime="00:02:32.85" />
                    <SPLIT distance="300" swimtime="00:03:51.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="442" reactiontime="+68" swimtime="00:01:08.32" resultid="17828" heatid="20093" lane="1" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4695538" athleteid="17740">
              <RESULTS>
                <RESULT eventid="3649" points="506" reactiontime="+65" swimtime="00:02:07.98" resultid="17741" heatid="19898" lane="8" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="521" reactiontime="+64" swimtime="00:04:33.36" resultid="17742" heatid="20057" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.99" />
                    <SPLIT distance="200" swimtime="00:02:13.38" />
                    <SPLIT distance="300" swimtime="00:03:24.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="458" reactiontime="+51" swimtime="00:05:16.31" resultid="17743" heatid="20118" lane="4" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="200" swimtime="00:02:36.51" />
                    <SPLIT distance="300" swimtime="00:04:07.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4938172" athleteid="17671">
              <RESULTS>
                <RESULT eventid="3628" points="228" reactiontime="+96" swimtime="00:01:35.83" resultid="17672" heatid="19866" lane="8" entrytime="00:01:35.12" />
                <RESULT eventid="3562" points="192" reactiontime="+82" swimtime="00:01:26.23" resultid="17673" heatid="19977" lane="7" entrytime="00:01:29.67" />
                <RESULT eventid="3578" points="338" reactiontime="+72" swimtime="00:05:15.85" resultid="17674" heatid="20055" lane="7" entrytime="00:05:26.86">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="200" swimtime="00:02:37.85" />
                    <SPLIT distance="300" swimtime="00:03:58.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="303" swimtime="00:06:02.94" resultid="17675" heatid="20116" lane="5" entrytime="00:06:20.79">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.24" />
                    <SPLIT distance="200" swimtime="00:02:55.89" />
                    <SPLIT distance="300" swimtime="00:04:42.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4843913" athleteid="17749">
              <RESULTS>
                <RESULT eventid="3628" points="404" reactiontime="+75" swimtime="00:01:19.18" resultid="17750" heatid="19870" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="3545" points="375" reactiontime="+70" swimtime="00:02:56.43" resultid="17751" heatid="19915" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="278" swimtime="00:01:19.49" resultid="17752" heatid="20014" lane="7" entrytime="00:01:32.91" />
                <RESULT eventid="3530" points="356" reactiontime="+75" swimtime="00:01:06.14" resultid="17753" heatid="20106" lane="8" entrytime="00:01:09.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4938673" athleteid="17810">
              <RESULTS>
                <RESULT eventid="3570" points="432" swimtime="00:02:29.34" resultid="17811" heatid="19882" lane="4" entrytime="00:02:30.51">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="480" swimtime="00:02:39.40" resultid="17812" heatid="19991" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="430" swimtime="00:01:16.95" resultid="17813" heatid="20010" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="3658" points="437" reactiontime="+62" swimtime="00:05:15.05" resultid="17814" heatid="20047" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.69" />
                    <SPLIT distance="200" swimtime="00:02:37.95" />
                    <SPLIT distance="300" swimtime="00:03:59.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4639374" athleteid="17563">
              <RESULTS>
                <RESULT eventid="3570" points="443" reactiontime="+72" swimtime="00:02:28.20" resultid="17564" heatid="19884" lane="8" entrytime="00:02:27.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="307" swimtime="00:01:23.09" resultid="17565" heatid="19971" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="3658" points="450" reactiontime="+68" swimtime="00:05:11.93" resultid="17566" heatid="20047" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.34" />
                    <SPLIT distance="200" swimtime="00:02:31.90" />
                    <SPLIT distance="300" swimtime="00:03:51.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="371" reactiontime="+68" swimtime="00:01:12.45" resultid="17567" heatid="20094" lane="8" entrytime="00:01:08.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4585059" athleteid="17788">
              <RESULTS>
                <RESULT eventid="3570" points="470" reactiontime="+75" swimtime="00:02:25.26" resultid="17789" heatid="19886" lane="2" entrytime="00:02:20.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="437" swimtime="00:02:44.37" resultid="17790" heatid="19991" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="484" swimtime="00:05:04.50" resultid="17791" heatid="20048" lane="5" entrytime="00:04:59.41">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                    <SPLIT distance="200" swimtime="00:02:30.69" />
                    <SPLIT distance="300" swimtime="00:03:48.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="446" swimtime="00:01:08.11" resultid="17792" heatid="20093" lane="4" entrytime="00:01:08.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4734887" athleteid="17581">
              <RESULTS>
                <RESULT eventid="3570" points="491" swimtime="00:02:23.16" resultid="17582" heatid="19885" lane="3" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="512" swimtime="00:02:35.96" resultid="17583" heatid="19992" lane="3" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="488" swimtime="00:01:13.79" resultid="17584" heatid="20011" lane="8" entrytime="00:01:13.00" />
                <RESULT eventid="3523" points="482" swimtime="00:01:06.41" resultid="17585" heatid="20097" lane="4" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4843896" athleteid="17815">
              <RESULTS>
                <RESULT eventid="3570" points="521" swimtime="00:02:20.34" resultid="17816" heatid="19886" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="467" swimtime="00:01:14.89" resultid="17817" heatid="20012" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="3586" points="407" reactiontime="+76" swimtime="00:02:44.24" resultid="17818" heatid="20064" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4810944" athleteid="17736">
              <RESULTS>
                <RESULT eventid="3649" points="418" reactiontime="+70" swimtime="00:02:16.32" resultid="17737" heatid="19896" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="365" swimtime="00:02:36.49" resultid="17738" heatid="19999" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                  </SPLITS>
                </RESULT>
                <RESULT comment=" - Wende mit einer Hand (Zeit: 15:18)" eventid="1081" reactiontime="+80" status="DSQ" swimtime="00:05:30.66" resultid="17739" heatid="20117" lane="7" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.01" />
                    <SPLIT distance="200" swimtime="00:02:40.40" />
                    <SPLIT distance="300" swimtime="00:04:16.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4695528" athleteid="17778">
              <RESULTS>
                <RESULT eventid="3621" points="436" reactiontime="+71" swimtime="00:01:24.95" resultid="17779" heatid="19860" lane="2" entrytime="00:01:27.75" />
                <RESULT eventid="3590" points="497" swimtime="00:00:29.95" resultid="17780" heatid="19934" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="3617" points="421" swimtime="00:00:33.43" resultid="17781" heatid="20029" lane="3" entrytime="00:00:32.97" />
                <RESULT eventid="3523" points="527" reactiontime="+68" swimtime="00:01:04.43" resultid="17782" heatid="20098" lane="8" entrytime="00:01:04.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" athleteid="17535">
              <RESULTS>
                <RESULT eventid="3628" points="162" swimtime="00:01:47.43" resultid="17536" heatid="19864" lane="4" entrytime="00:01:42.57" />
                <RESULT eventid="3594" points="233" swimtime="00:00:33.97" resultid="17537" heatid="19949" lane="5" entrytime="00:00:34.82" />
                <RESULT eventid="3530" points="241" swimtime="00:01:15.33" resultid="17538" heatid="20104" lane="8" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4809423" athleteid="17553">
              <RESULTS>
                <RESULT eventid="3570" points="597" reactiontime="+80" swimtime="00:02:14.11" resultid="17554" heatid="19888" lane="2" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="459" reactiontime="+83" swimtime="00:01:12.67" resultid="17555" heatid="19973" lane="6" entrytime="00:01:12.50" />
                <RESULT eventid="3658" points="623" reactiontime="+66" swimtime="00:04:39.95" resultid="17556" heatid="20050" lane="3" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="200" swimtime="00:02:16.41" />
                    <SPLIT distance="300" swimtime="00:03:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" points="383" reactiontime="+76" swimtime="00:02:47.63" resultid="17557" heatid="20065" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4809375" athleteid="17641">
              <RESULTS>
                <RESULT eventid="9711" points="345" reactiontime="+66" swimtime="00:02:42.40" resultid="17642" heatid="19828" lane="1" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="310" reactiontime="+57" swimtime="00:01:26.49" resultid="17643" heatid="19868" lane="2" entrytime="00:01:25.50" />
                <RESULT eventid="3562" points="339" reactiontime="+61" swimtime="00:01:11.41" resultid="17644" heatid="19979" lane="4" entrytime="00:01:08.00" />
                <RESULT eventid="3613" points="373" swimtime="00:00:31.14" resultid="17645" heatid="20037" lane="8" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5001366" athleteid="17503">
              <RESULTS>
                <RESULT eventid="3621" points="242" swimtime="00:01:43.38" resultid="17504" heatid="19857" lane="8" entrytime="00:01:37.80" />
                <RESULT eventid="3570" points="264" reactiontime="+87" swimtime="00:02:55.96" resultid="17505" heatid="19879" lane="6" entrytime="00:02:50.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="294" reactiontime="+68" swimtime="00:01:18.30" resultid="17506" heatid="20089" lane="2" entrytime="00:01:15.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4907136" athleteid="17568">
              <RESULTS>
                <RESULT eventid="3570" points="392" reactiontime="+60" swimtime="00:02:34.26" resultid="17569" heatid="19881" lane="1" entrytime="00:02:40.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="361" swimtime="00:00:33.31" resultid="17570" heatid="19927" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="3505" points="407" swimtime="00:02:48.29" resultid="17571" heatid="19988" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="422" swimtime="00:01:17.44" resultid="17572" heatid="20008" lane="1" entrytime="00:01:22.65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5001364" athleteid="17523">
              <RESULTS>
                <RESULT eventid="3621" points="240" reactiontime="+98" swimtime="00:01:43.61" resultid="17524" heatid="19856" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="3590" points="269" swimtime="00:00:36.76" resultid="17525" heatid="19924" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="3514" points="266" swimtime="00:00:46.32" resultid="17526" heatid="20071" lane="2" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4585067" athleteid="17716">
              <RESULTS>
                <RESULT eventid="3628" points="437" reactiontime="+63" swimtime="00:01:17.17" resultid="17717" heatid="19870" lane="8" entrytime="00:01:20.00" />
                <RESULT eventid="3545" points="449" reactiontime="+72" swimtime="00:02:46.24" resultid="17718" heatid="19914" lane="4" entrytime="00:02:53.48">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="324" swimtime="00:01:15.59" resultid="17719" heatid="20018" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="3588" points="375" reactiontime="+55" swimtime="00:02:34.51" resultid="17720" heatid="20066" lane="4" entrytime="00:02:38.09">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4489640" athleteid="17676">
              <RESULTS>
                <RESULT eventid="3628" points="405" reactiontime="+52" swimtime="00:01:19.15" resultid="17677" heatid="19871" lane="4" entrytime="00:01:14.00" />
                <RESULT eventid="3594" points="459" swimtime="00:00:27.09" resultid="17678" heatid="19958" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="3613" points="480" swimtime="00:00:28.64" resultid="17679" heatid="20039" lane="8" entrytime="00:00:27.45" />
                <RESULT eventid="3530" points="491" reactiontime="+71" swimtime="00:00:59.45" resultid="17680" heatid="20111" lane="7" entrytime="00:00:56.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4489647" athleteid="17681">
              <RESULTS>
                <RESULT eventid="9711" points="387" swimtime="00:02:36.43" resultid="17682" heatid="19829" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="366" reactiontime="+69" swimtime="00:01:21.86" resultid="17683" heatid="19870" lane="7" entrytime="00:01:20.00" />
                <RESULT eventid="3605" points="394" swimtime="00:01:10.82" resultid="17684" heatid="20020" lane="2" entrytime="00:01:11.00" />
                <RESULT eventid="3530" points="431" reactiontime="+52" swimtime="00:01:02.07" resultid="17685" heatid="20108" lane="3" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4760057" athleteid="17611">
              <RESULTS>
                <RESULT eventid="9711" points="427" reactiontime="+76" swimtime="00:02:31.35" resultid="17612" heatid="19830" lane="8" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="478" swimtime="00:00:26.73" resultid="17613" heatid="19956" lane="4" entrytime="00:00:26.50" />
                <RESULT eventid="3613" points="414" swimtime="00:00:30.08" resultid="17614" heatid="20037" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="3530" points="516" reactiontime="+74" swimtime="00:00:58.47" resultid="17615" heatid="20110" lane="5" entrytime="00:00:57.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4500966" athleteid="17686">
              <RESULTS>
                <RESULT eventid="3649" points="564" reactiontime="+62" swimtime="00:02:03.39" resultid="17687" heatid="19898" lane="3" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="517" swimtime="00:02:19.38" resultid="17688" heatid="20001" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="513" swimtime="00:01:04.85" resultid="17689" heatid="20022" lane="8" entrytime="00:01:04.00" />
                <RESULT eventid="3519" points="529" swimtime="00:00:32.96" resultid="17690" heatid="20084" lane="1" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5006990" athleteid="17651">
              <RESULTS>
                <RESULT eventid="3570" points="339" swimtime="00:02:41.89" resultid="17652" heatid="19879" lane="3" entrytime="00:02:50.64">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="330" swimtime="00:01:21.09" resultid="17653" heatid="19970" lane="1" entrytime="00:01:28.81" />
                <RESULT eventid="3598" points="333" swimtime="00:01:23.78" resultid="17654" heatid="20006" lane="3" entrytime="00:01:25.19" />
                <RESULT eventid="3636" points="358" reactiontime="+75" swimtime="00:06:19.28" resultid="17655" heatid="20114" lane="1" entrytime="00:06:13.51">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.73" />
                    <SPLIT distance="200" swimtime="00:03:04.11" />
                    <SPLIT distance="300" swimtime="00:04:51.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5039264" athleteid="17806">
              <RESULTS>
                <RESULT eventid="3570" points="405" swimtime="00:02:32.69" resultid="17807" heatid="19884" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="382" swimtime="00:02:51.87" resultid="17808" heatid="19990" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" status="DNS" swimtime="00:00:00.00" resultid="17809" heatid="20046" lane="7" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4495032" athleteid="17548">
              <RESULTS>
                <RESULT eventid="3570" points="518" reactiontime="+65" swimtime="00:02:20.63" resultid="17549" heatid="19887" lane="1" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="440" swimtime="00:02:44.05" resultid="17550" heatid="19992" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" status="DNS" swimtime="00:00:00.00" resultid="17551" heatid="20012" lane="5" entrytime="00:01:09.50" />
                <RESULT eventid="3523" points="544" reactiontime="+75" swimtime="00:01:03.78" resultid="17552" heatid="20099" lane="8" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4844648" athleteid="17596">
              <RESULTS>
                <RESULT eventid="9711" points="411" swimtime="00:02:33.29" resultid="17597" heatid="19829" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="365" reactiontime="+78" swimtime="00:01:09.65" resultid="17598" heatid="19979" lane="7" entrytime="00:01:09.00" />
                <RESULT eventid="3605" points="391" swimtime="00:01:11.01" resultid="17599" heatid="20019" lane="5" entrytime="00:01:12.00" />
                <RESULT eventid="1081" points="416" reactiontime="+76" swimtime="00:05:26.41" resultid="17600" heatid="20118" lane="2" entrytime="00:05:19.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                    <SPLIT distance="200" swimtime="00:02:37.93" />
                    <SPLIT distance="300" swimtime="00:04:13.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4500994" athleteid="17773">
              <RESULTS>
                <RESULT eventid="3639" points="420" reactiontime="+66" swimtime="00:02:48.35" resultid="17774" heatid="19819" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="507" swimtime="00:02:36.44" resultid="17775" heatid="19993" lane="8" entrytime="00:02:32.44">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="476" swimtime="00:01:14.41" resultid="17776" heatid="20011" lane="3" entrytime="00:01:11.79" />
                <RESULT eventid="3636" points="440" reactiontime="+49" swimtime="00:05:54.14" resultid="17777" heatid="20115" lane="1" entrytime="00:05:39.55">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.80" />
                    <SPLIT distance="200" swimtime="00:02:48.10" />
                    <SPLIT distance="300" swimtime="00:04:34.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4695532" athleteid="17793">
              <RESULTS>
                <RESULT eventid="3547" points="612" swimtime="00:00:31.86" resultid="17794" heatid="19844" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="3590" points="529" swimtime="00:00:29.33" resultid="17795" heatid="19933" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="3658" points="624" reactiontime="+74" swimtime="00:04:39.76" resultid="17796" heatid="20050" lane="6" entrytime="00:04:41.72">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.34" />
                    <SPLIT distance="200" swimtime="00:02:17.05" />
                    <SPLIT distance="300" swimtime="00:03:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" points="594" swimtime="00:02:24.89" resultid="17797" heatid="20065" lane="5" entrytime="00:02:21.51">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4929333" athleteid="17636">
              <RESULTS>
                <RESULT eventid="3649" points="422" reactiontime="+76" swimtime="00:02:15.90" resultid="17637" heatid="19897" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="403" swimtime="00:00:28.29" resultid="17638" heatid="19955" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="3578" points="457" reactiontime="+78" swimtime="00:04:45.51" resultid="17639" heatid="20056" lane="6" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="200" swimtime="00:02:20.39" />
                    <SPLIT distance="300" swimtime="00:03:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3588" points="313" swimtime="00:02:44.19" resultid="17640" heatid="20067" lane="2" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="5001068" athleteid="17539">
              <RESULTS>
                <RESULT eventid="3551" points="179" swimtime="00:00:42.59" resultid="17540" heatid="19847" lane="6" entrytime="00:00:42.40" />
                <RESULT eventid="3605" points="197" swimtime="00:01:29.20" resultid="17541" heatid="20016" lane="8" entrytime="00:01:25.80" />
                <RESULT eventid="3530" points="255" swimtime="00:01:13.94" resultid="17542" heatid="20102" lane="2" entrytime="00:01:19.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="5001070" athleteid="17531">
              <RESULTS>
                <RESULT eventid="3628" points="398" reactiontime="+72" swimtime="00:01:19.62" resultid="17532" heatid="19871" lane="1" entrytime="00:01:18.00" />
                <RESULT eventid="3594" points="392" swimtime="00:00:28.55" resultid="17533" heatid="19953" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="3519" points="469" swimtime="00:00:34.31" resultid="17534" heatid="20083" lane="4" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4735391" athleteid="17573">
              <RESULTS>
                <RESULT eventid="3570" points="468" reactiontime="+67" swimtime="00:02:25.49" resultid="17574" heatid="19884" lane="3" entrytime="00:02:25.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="393" reactiontime="+71" swimtime="00:01:16.51" resultid="17575" heatid="19972" lane="6" entrytime="00:01:16.66" />
                <RESULT eventid="3617" points="437" swimtime="00:00:33.02" resultid="17576" heatid="20029" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="3523" points="462" reactiontime="+80" swimtime="00:01:07.32" resultid="17577" heatid="20095" lane="6" entrytime="00:01:07.60" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="12820" points="584" swimtime="00:04:07.88" resultid="19692" heatid="20141" lane="5" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="200" swimtime="00:02:10.43" />
                    <SPLIT distance="300" swimtime="00:03:10.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17706" number="1" />
                    <RELAYPOSITION athleteid="17691" number="2" reactiontime="+11" />
                    <RELAYPOSITION athleteid="17763" number="3" />
                    <RELAYPOSITION athleteid="17626" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12864" points="572" reactiontime="+63" swimtime="00:03:46.76" resultid="19700" heatid="20137" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.87" />
                    <SPLIT distance="200" swimtime="00:01:52.11" />
                    <SPLIT distance="300" swimtime="00:02:49.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17686" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="17701" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="17626" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="17696" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="12820" points="528" swimtime="00:04:16.37" resultid="19693" heatid="20141" lane="3" entrytime="00:04:09.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.63" />
                    <SPLIT distance="200" swimtime="00:02:15.15" />
                    <SPLIT distance="300" swimtime="00:03:18.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17686" number="1" />
                    <RELAYPOSITION athleteid="17701" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="17696" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="17611" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12864" points="494" reactiontime="+48" swimtime="00:03:58.10" resultid="19701" heatid="20137" lane="2" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.48" />
                    <SPLIT distance="200" swimtime="00:01:58.06" />
                    <SPLIT distance="300" swimtime="00:02:58.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17763" number="1" reactiontime="+48" />
                    <RELAYPOSITION athleteid="17681" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="17596" number="3" reactiontime="-1" />
                    <RELAYPOSITION athleteid="17676" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="12820" points="338" swimtime="00:04:57.41" resultid="19695" heatid="20140" lane="5" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.88" />
                    <SPLIT distance="200" swimtime="00:02:34.28" />
                    <SPLIT distance="300" swimtime="00:03:48.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17527" number="1" />
                    <RELAYPOSITION athleteid="17531" number="2" />
                    <RELAYPOSITION athleteid="17519" number="3" />
                    <RELAYPOSITION athleteid="17586" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12864" points="344" reactiontime="+63" swimtime="00:04:28.52" resultid="19703" heatid="20136" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="200" swimtime="00:02:15.15" />
                    <SPLIT distance="300" swimtime="00:03:25.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17527" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="17666" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="17671" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="17531" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="12820" points="444" swimtime="00:04:31.68" resultid="19694" heatid="20141" lane="1" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.97" />
                    <SPLIT distance="200" swimtime="00:02:27.06" />
                    <SPLIT distance="300" swimtime="00:03:30.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17726" number="1" />
                    <RELAYPOSITION athleteid="17749" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="17721" number="3" reactiontime="+7" />
                    <RELAYPOSITION athleteid="17636" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12864" points="485" reactiontime="+48" swimtime="00:03:59.43" resultid="19702" heatid="20137" lane="7" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.27" />
                    <SPLIT distance="200" swimtime="00:01:57.72" />
                    <SPLIT distance="300" swimtime="00:02:58.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17740" number="1" reactiontime="+48" />
                    <RELAYPOSITION athleteid="17611" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="17711" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="17758" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="3574" points="585" swimtime="00:04:37.48" resultid="19696" heatid="20139" lane="4" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.51" />
                    <SPLIT distance="200" swimtime="00:02:28.81" />
                    <SPLIT distance="300" swimtime="00:03:35.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17793" number="1" />
                    <RELAYPOSITION athleteid="17558" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="17845" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="17553" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12862" points="629" swimtime="00:04:07.05" resultid="19704" heatid="20135" lane="4" entrytime="00:04:06.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.44" />
                    <SPLIT distance="200" swimtime="00:02:05.24" />
                    <SPLIT distance="300" swimtime="00:03:05.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17793" number="1" />
                    <RELAYPOSITION athleteid="17553" number="2" />
                    <RELAYPOSITION athleteid="17845" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="17558" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="3574" points="449" swimtime="00:05:03.19" resultid="19697" heatid="20139" lane="8" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="200" swimtime="00:02:37.96" />
                    <SPLIT distance="300" swimtime="00:03:58.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17543" number="1" />
                    <RELAYPOSITION athleteid="17778" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="17783" number="3" reactiontime="-3" />
                    <RELAYPOSITION athleteid="17548" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12862" points="473" reactiontime="+50" swimtime="00:04:31.67" resultid="19705" heatid="20135" lane="2" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.76" />
                    <SPLIT distance="200" swimtime="00:02:16.60" />
                    <SPLIT distance="300" swimtime="00:03:26.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17773" number="1" reactiontime="+50" />
                    <RELAYPOSITION athleteid="17788" number="2" />
                    <RELAYPOSITION athleteid="17563" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="17768" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="3574" points="493" swimtime="00:04:53.88" resultid="19698" heatid="20138" lane="5" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.12" />
                    <SPLIT distance="200" swimtime="00:02:35.91" />
                    <SPLIT distance="300" swimtime="00:03:47.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17581" number="1" />
                    <RELAYPOSITION athleteid="17798" number="2" />
                    <RELAYPOSITION athleteid="17815" number="3" />
                    <RELAYPOSITION athleteid="17573" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12862" points="334" swimtime="00:05:04.96" resultid="19707" heatid="20134" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="200" swimtime="00:02:31.59" />
                    <SPLIT distance="300" swimtime="00:03:46.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17841" number="1" />
                    <RELAYPOSITION athleteid="17503" number="2" />
                    <RELAYPOSITION athleteid="17651" number="3" />
                    <RELAYPOSITION athleteid="17646" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="3574" points="389" swimtime="00:05:17.98" resultid="19699" heatid="20138" lane="2" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="200" swimtime="00:02:46.04" />
                    <SPLIT distance="300" swimtime="00:04:04.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17837" number="1" />
                    <RELAYPOSITION athleteid="17829" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="17507" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="17833" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12862" points="457" reactiontime="+58" swimtime="00:04:34.69" resultid="19706" heatid="20135" lane="8" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="200" swimtime="00:02:20.42" />
                    <SPLIT distance="300" swimtime="00:03:27.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17810" number="1" reactiontime="+58" />
                    <RELAYPOSITION athleteid="17591" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="17581" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="17824" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="BREGENZ" nation="AUT" region="VLSV" clubid="13981" swrid="66431" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2000-10-04" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="4520432" athleteid="17276">
              <RESULTS>
                <RESULT eventid="3639" points="362" reactiontime="+55" swimtime="00:02:56.91" resultid="17277" heatid="19814" lane="8" entrytime="00:03:03.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="407" reactiontime="+53" swimtime="00:01:26.92" resultid="17278" heatid="19859" lane="1" entrytime="00:01:31.49" entrycourse="LCM" />
                <RESULT eventid="3538" points="402" reactiontime="+69" swimtime="00:03:09.80" resultid="17279" heatid="19907" lane="6" entrytime="00:03:16.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="395" swimtime="00:00:32.34" resultid="17280" heatid="19927" lane="4" entrytime="00:00:33.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-09-03" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="4746948" athleteid="17243">
              <RESULTS>
                <RESULT eventid="9711" points="296" reactiontime="+68" swimtime="00:02:50.88" resultid="17244" heatid="19825" lane="4" entrytime="00:03:02.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="246" swimtime="00:00:38.32" resultid="17245" heatid="19848" lane="7" entrytime="00:00:40.11" entrycourse="LCM" />
                <RESULT eventid="3649" points="309" reactiontime="+74" swimtime="00:02:30.76" resultid="17246" heatid="19893" lane="8" entrytime="00:02:37.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="293" swimtime="00:00:31.45" resultid="17247" heatid="19951" lane="7" entrytime="00:00:32.03" entrycourse="LCM" />
                <RESULT eventid="3512" points="240" swimtime="00:02:59.85" resultid="17248" heatid="19996" lane="8" entrytime="00:03:09.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="5172648" athleteid="17254">
              <RESULTS>
                <RESULT eventid="3621" points="239" reactiontime="+83" swimtime="00:01:43.75" resultid="17255" heatid="19855" lane="7" entrytime="00:01:42.99" entrycourse="SCM" />
                <RESULT eventid="3570" points="258" reactiontime="+87" swimtime="00:02:57.44" resultid="17256" heatid="19880" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="402" swimtime="00:00:32.15" resultid="17257" heatid="19927" lane="5" entrytime="00:00:33.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-05-15" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="4769224" athleteid="17249">
              <RESULTS>
                <RESULT eventid="9711" points="499" reactiontime="+70" swimtime="00:02:23.67" resultid="17250" heatid="19831" lane="2" entrytime="00:02:24.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="500" reactiontime="+75" swimtime="00:01:13.80" resultid="17251" heatid="19872" lane="8" entrytime="00:01:13.09" entrycourse="LCM" />
                <RESULT eventid="3545" points="451" reactiontime="+72" swimtime="00:02:45.93" resultid="17252" heatid="19915" lane="5" entrytime="00:02:46.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="398" reactiontime="+75" swimtime="00:01:07.68" resultid="17253" heatid="19978" lane="3" entrytime="00:01:11.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-28" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="4557331" athleteid="17258">
              <RESULTS>
                <RESULT eventid="3551" points="401" swimtime="00:00:32.59" resultid="17259" heatid="19851" lane="1" entrytime="00:00:31.30" entrycourse="SCM" />
                <RESULT eventid="3649" points="378" reactiontime="+61" swimtime="00:02:21.01" resultid="17260" heatid="19895" lane="4" entrytime="00:02:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="414" swimtime="00:00:28.04" resultid="17261" heatid="19956" lane="6" entrytime="00:00:27.14" entrycourse="SCM" />
                <RESULT eventid="3512" points="329" swimtime="00:02:42.00" resultid="17262" heatid="20000" lane="8" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-02-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="4769221" athleteid="17263">
              <RESULTS>
                <RESULT eventid="3639" points="421" reactiontime="+58" swimtime="00:02:48.24" resultid="17264" heatid="19816" lane="4" entrytime="00:02:52.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="435" swimtime="00:00:35.70" resultid="17265" heatid="19842" lane="3" entrytime="00:00:35.57" entrycourse="LCM" />
                <RESULT eventid="3505" points="493" swimtime="00:02:37.96" resultid="17266" heatid="19991" lane="5" entrytime="00:02:38.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="461" swimtime="00:01:15.21" resultid="17267" heatid="20010" lane="7" entrytime="00:01:15.91" entrycourse="LCM" />
                <RESULT eventid="3617" points="402" swimtime="00:00:33.95" resultid="17268" heatid="20027" lane="4" entrytime="00:00:36.30" entrycourse="LCM" />
                <RESULT eventid="3523" points="458" reactiontime="+69" swimtime="00:01:07.51" resultid="17269" heatid="20094" lane="2" entrytime="00:01:08.44" entrycourse="LCM" />
                <RESULT eventid="3636" points="440" reactiontime="+57" swimtime="00:05:54.11" resultid="17270" heatid="20114" lane="7" entrytime="00:06:04.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.46" />
                    <SPLIT distance="200" swimtime="00:02:50.51" />
                    <SPLIT distance="300" swimtime="00:04:38.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="5127529" athleteid="17271">
              <RESULTS>
                <RESULT eventid="3639" points="288" reactiontime="+77" swimtime="00:03:10.98" resultid="17272" heatid="19810" lane="8" entrytime="00:03:28.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="298" swimtime="00:01:36.48" resultid="17273" heatid="19855" lane="2" entrytime="00:01:42.91" entrycourse="LCM" />
                <RESULT eventid="3538" points="321" reactiontime="+70" swimtime="00:03:24.45" resultid="17274" heatid="19905" lane="2" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="322" swimtime="00:00:34.60" resultid="17275" heatid="19923" lane="4" entrytime="00:00:37.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCSH" nation="SUI" region="ROS" clubid="14333" swrid="65668" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2004-08-04" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4894102" athleteid="18253">
              <RESULTS>
                <RESULT eventid="3551" points="227" swimtime="00:00:39.38" resultid="18254" heatid="19847" lane="5" entrytime="00:00:42.07" />
                <RESULT eventid="3649" points="247" swimtime="00:02:42.45" resultid="18255" heatid="19890" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="200" reactiontime="+70" swimtime="00:03:37.55" resultid="18256" heatid="19911" lane="5" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="230" swimtime="00:03:02.51" resultid="18257" heatid="19997" lane="7" entrytime="00:02:58.02">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="224" swimtime="00:01:25.49" resultid="18258" heatid="20015" lane="4" entrytime="00:01:25.82" />
                <RESULT eventid="3578" points="265" reactiontime="+69" swimtime="00:05:42.23" resultid="18259" heatid="20054" lane="7" entrytime="00:05:39.38">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.75" />
                    <SPLIT distance="200" swimtime="00:02:48.50" />
                    <SPLIT distance="300" swimtime="00:04:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="173" swimtime="00:00:47.81" resultid="18260" heatid="20078" lane="4" entrytime="00:00:50.13" />
                <RESULT eventid="3530" points="239" swimtime="00:01:15.51" resultid="18261" heatid="20103" lane="3" entrytime="00:01:15.62" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="4968038" athleteid="18220">
              <RESULTS>
                <RESULT eventid="3639" points="231" swimtime="00:03:25.42" resultid="18221" heatid="19810" lane="4" entrytime="00:03:18.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="291" reactiontime="+77" swimtime="00:02:50.46" resultid="18222" heatid="19878" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="264" swimtime="00:00:36.97" resultid="18223" heatid="19922" lane="4" entrytime="00:00:39.04" />
                <RESULT eventid="3505" points="255" swimtime="00:03:16.74" resultid="18224" heatid="19983" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="234" swimtime="00:01:34.27" resultid="18225" heatid="20003" lane="3" entrytime="00:01:34.52" />
                <RESULT eventid="3658" points="308" swimtime="00:05:54.03" resultid="18226" heatid="20041" lane="3" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="200" swimtime="00:02:54.52" />
                    <SPLIT distance="300" swimtime="00:04:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="223" swimtime="00:00:49.11" resultid="18227" heatid="20070" lane="1" entrytime="00:00:52.34" />
                <RESULT eventid="3523" points="278" reactiontime="+75" swimtime="00:01:19.77" resultid="18228" heatid="20087" lane="5" entrytime="00:01:20.19" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-11-18" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="5133828" athleteid="18440">
              <RESULTS>
                <RESULT eventid="9711" points="167" swimtime="00:03:26.84" resultid="18441" heatid="19824" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="230" swimtime="00:02:46.38" resultid="18442" heatid="19890" lane="6" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="217" swimtime="00:00:34.76" resultid="18443" heatid="19949" lane="4" entrytime="00:00:34.79" />
                <RESULT eventid="3562" points="86" swimtime="00:01:52.50" resultid="18444" heatid="19976" lane="4" entrytime="00:01:40.00" />
                <RESULT eventid="3613" points="138" swimtime="00:00:43.38" resultid="18445" heatid="20034" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="3578" points="241" swimtime="00:05:53.42" resultid="18446" heatid="20052" lane="7" entrytime="00:06:02.64">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.78" />
                    <SPLIT distance="200" swimtime="00:02:55.61" />
                    <SPLIT distance="300" swimtime="00:04:26.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="131" swimtime="00:00:52.39" resultid="18447" heatid="20077" lane="4" entrytime="00:00:52.72" />
                <RESULT eventid="3530" points="209" swimtime="00:01:18.93" resultid="18448" heatid="20102" lane="3" entrytime="00:01:18.56" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-12-11" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="26699" swrid="4465306" athleteid="18262">
              <RESULTS>
                <RESULT eventid="3547" points="478" swimtime="00:00:34.60" resultid="18263" heatid="19843" lane="1" entrytime="00:00:34.72" entrycourse="LCM" />
                <RESULT eventid="3570" points="553" reactiontime="+83" swimtime="00:02:17.61" resultid="18264" heatid="19886" lane="6" entrytime="00:02:20.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="476" swimtime="00:00:30.38" resultid="18265" heatid="19932" lane="6" entrytime="00:00:30.73" entrycourse="LCM" />
                <RESULT eventid="3505" points="566" swimtime="00:02:30.85" resultid="18266" heatid="19992" lane="8" entrytime="00:02:36.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="510" swimtime="00:01:12.73" resultid="18267" heatid="20011" lane="2" entrytime="00:01:12.46" entrycourse="LCM" />
                <RESULT eventid="3658" points="559" reactiontime="+83" swimtime="00:04:50.30" resultid="18268" heatid="20049" lane="6" entrytime="00:04:51.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.55" />
                    <SPLIT distance="200" swimtime="00:02:21.66" />
                    <SPLIT distance="300" swimtime="00:03:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="415" swimtime="00:00:39.95" resultid="18269" heatid="20072" lane="3" entrytime="00:00:43.24" />
                <RESULT eventid="3523" points="504" reactiontime="+77" swimtime="00:01:05.40" resultid="18270" heatid="20096" lane="6" entrytime="00:01:06.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-08-28" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="5003011" athleteid="18431">
              <RESULTS>
                <RESULT eventid="9711" points="208" swimtime="00:03:12.34" resultid="18432" heatid="19825" lane="8" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="275" swimtime="00:02:36.74" resultid="18433" heatid="19891" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="215" swimtime="00:00:34.90" resultid="18434" heatid="19949" lane="1" entrytime="00:00:35.22" />
                <RESULT eventid="3512" points="215" swimtime="00:03:06.67" resultid="18435" heatid="19996" lane="1" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="200" swimtime="00:01:28.76" resultid="18436" heatid="20015" lane="1" entrytime="00:01:29.38" />
                <RESULT eventid="3578" points="303" swimtime="00:05:27.57" resultid="18437" heatid="20054" lane="6" entrytime="00:05:33.57">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="200" swimtime="00:02:43.06" />
                    <SPLIT distance="300" swimtime="00:04:07.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="157" swimtime="00:00:49.39" resultid="18438" heatid="20079" lane="1" entrytime="00:00:48.64" />
                <RESULT eventid="3530" points="251" swimtime="00:01:14.27" resultid="18439" heatid="20103" lane="4" entrytime="00:01:15.06" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-31" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="24812" swrid="4354800" athleteid="18318">
              <RESULTS>
                <RESULT eventid="3639" points="511" reactiontime="+61" swimtime="00:02:37.79" resultid="18319" heatid="19821" lane="3" entrytime="00:02:35.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="532" reactiontime="+76" swimtime="00:02:19.42" resultid="18320" heatid="19887" lane="7" entrytime="00:02:16.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="517" swimtime="00:00:29.55" resultid="18321" heatid="19937" lane="8" entrytime="00:00:29.39" entrycourse="LCM" />
                <RESULT eventid="3555" points="462" reactiontime="+74" swimtime="00:01:12.49" resultid="18322" heatid="19974" lane="2" entrytime="00:01:10.00" entrycourse="LCM" />
                <RESULT eventid="3598" points="399" swimtime="00:01:18.91" resultid="18323" heatid="20010" lane="3" entrytime="00:01:14.81" />
                <RESULT eventid="3658" status="DNS" swimtime="00:00:00.00" resultid="18324" heatid="20050" lane="8" entrytime="00:04:47.59" entrycourse="LCM" />
                <RESULT eventid="3586" status="DNS" swimtime="00:00:00.00" resultid="18325" heatid="20065" lane="3" entrytime="00:02:34.03" entrycourse="LCM" />
                <RESULT eventid="3523" status="DNS" swimtime="00:00:00.00" resultid="18326" heatid="20098" lane="6" entrytime="00:01:03.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-04-17" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="13475" swrid="4022292" athleteid="18391">
              <RESULTS>
                <RESULT eventid="3639" points="706" swimtime="00:02:21.67" resultid="18392" heatid="19822" lane="5" entrytime="00:02:20.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="613" swimtime="00:01:15.83" resultid="18393" heatid="19863" lane="4" entrytime="00:01:14.09" entrycourse="LCM" />
                <RESULT eventid="3538" points="659" swimtime="00:02:41.00" resultid="18394" heatid="19910" lane="4" entrytime="00:02:42.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="621" swimtime="00:00:27.80" resultid="18395" heatid="19935" lane="4" entrytime="00:00:27.18" entrycourse="LCM" />
                <RESULT eventid="3555" points="632" reactiontime="+58" swimtime="00:01:05.30" resultid="18396" heatid="19975" lane="3" entrytime="00:01:04.55" entrycourse="LCM" />
                <RESULT eventid="3658" points="699" reactiontime="+57" swimtime="00:04:29.45" resultid="18397" heatid="20050" lane="4" entrytime="00:04:23.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.20" />
                    <SPLIT distance="200" swimtime="00:02:12.71" />
                    <SPLIT distance="300" swimtime="00:03:21.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" points="623" reactiontime="+57" swimtime="00:02:22.61" resultid="18398" heatid="20065" lane="4" entrytime="00:02:19.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3636" points="713" reactiontime="+72" swimtime="00:05:01.55" resultid="18399" heatid="20115" lane="4" entrytime="00:04:55.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="200" swimtime="00:02:26.48" />
                    <SPLIT distance="300" swimtime="00:03:53.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15921" points="614" swimtime="00:00:27.91" resultid="20166" heatid="20120" lane="3" late="yes" />
                <RESULT eventid="15972" points="553" swimtime="00:00:28.91" resultid="20167" heatid="20122" lane="3" late="yes" />
                <RESULT eventid="15975" points="579" swimtime="00:00:28.47" resultid="20168" heatid="20124" lane="3" late="yes" />
                <RESULT eventid="15978" points="599" swimtime="00:00:28.14" resultid="20169" heatid="20126" lane="3" late="yes" />
                <RESULT eventid="15981" points="613" swimtime="00:00:27.92" resultid="20170" heatid="20128" lane="3" late="yes" />
                <RESULT eventid="15984" points="617" swimtime="00:00:27.87" resultid="20171" heatid="20130" lane="3" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-26" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="28176" swrid="4688318" athleteid="18288">
              <RESULTS>
                <RESULT eventid="3639" points="461" reactiontime="+61" swimtime="00:02:43.30" resultid="18289" heatid="19820" lane="1" entrytime="00:02:38.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="502" reactiontime="+57" swimtime="00:01:21.08" resultid="18290" heatid="19863" lane="7" entrytime="00:01:18.56" entrycourse="SCM" />
                <RESULT eventid="3538" points="491" swimtime="00:02:57.61" resultid="18291" heatid="19910" lane="3" entrytime="00:02:47.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="354" swimtime="00:01:19.22" resultid="18292" heatid="19972" lane="3" entrytime="00:01:16.42" entrycourse="LCM" />
                <RESULT eventid="3658" points="495" reactiontime="+57" swimtime="00:05:02.30" resultid="18293" heatid="20049" lane="8" entrytime="00:04:58.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="200" swimtime="00:02:26.86" />
                    <SPLIT distance="300" swimtime="00:03:44.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="534" swimtime="00:00:36.71" resultid="18294" heatid="20075" lane="3" entrytime="00:00:36.70" entrycourse="LCM" />
                <RESULT eventid="3523" points="487" reactiontime="+60" swimtime="00:01:06.14" resultid="18295" heatid="20097" lane="3" entrytime="00:01:05.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-06-29" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="27618" swrid="4621600" athleteid="18400">
              <RESULTS>
                <RESULT eventid="3639" points="606" reactiontime="+86" swimtime="00:02:29.04" resultid="18401" heatid="19822" lane="6" entrytime="00:02:29.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="578" swimtime="00:01:17.33" resultid="18402" heatid="19863" lane="5" entrytime="00:01:15.22" entrycourse="LCM" />
                <RESULT eventid="3538" points="607" swimtime="00:02:45.46" resultid="18403" heatid="19910" lane="5" entrytime="00:02:42.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="527" swimtime="00:00:29.36" resultid="18404" heatid="19936" lane="1" entrytime="00:00:29.22" entrycourse="LCM" />
                <RESULT eventid="3617" points="486" swimtime="00:00:31.87" resultid="18405" heatid="20030" lane="2" entrytime="00:00:31.68" entrycourse="LCM" />
                <RESULT eventid="3658" points="536" reactiontime="+80" swimtime="00:04:54.25" resultid="18406" heatid="20049" lane="5" entrytime="00:04:49.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="200" swimtime="00:02:24.08" />
                    <SPLIT distance="300" swimtime="00:03:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="605" swimtime="00:00:35.22" resultid="18407" heatid="20075" lane="5" entrytime="00:00:35.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-12-16" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="4894108" athleteid="18345">
              <RESULTS>
                <RESULT eventid="3639" points="479" reactiontime="+68" swimtime="00:02:41.19" resultid="18346" heatid="19820" lane="8" entrytime="00:02:38.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="495" swimtime="00:02:22.77" resultid="18347" heatid="19886" lane="4" entrytime="00:02:17.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="497" swimtime="00:00:29.94" resultid="18348" heatid="19935" lane="2" entrytime="00:00:28.86" entrycourse="SCM" />
                <RESULT eventid="3555" points="372" reactiontime="+65" swimtime="00:01:17.94" resultid="18349" heatid="19973" lane="4" entrytime="00:01:11.35" entrycourse="LCM" />
                <RESULT eventid="3598" points="450" swimtime="00:01:15.80" resultid="18350" heatid="20010" lane="5" entrytime="00:01:14.40" entrycourse="LCM" />
                <RESULT eventid="3658" points="520" swimtime="00:04:57.33" resultid="18351" heatid="20049" lane="3" entrytime="00:04:50.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.17" />
                    <SPLIT distance="200" swimtime="00:02:28.02" />
                    <SPLIT distance="300" swimtime="00:03:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="531" reactiontime="+71" swimtime="00:01:04.29" resultid="18352" heatid="20099" lane="7" entrytime="00:01:02.80" entrycourse="LCM" />
                <RESULT eventid="3636" points="454" reactiontime="+77" swimtime="00:05:50.46" resultid="18353" heatid="20115" lane="7" entrytime="00:05:39.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                    <SPLIT distance="200" swimtime="00:02:52.85" />
                    <SPLIT distance="300" swimtime="00:04:36.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-07-28" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="23350" swrid="4228679" athleteid="18104">
              <RESULTS>
                <RESULT eventid="3639" points="429" reactiontime="+63" swimtime="00:02:47.26" resultid="18105" heatid="19821" lane="2" entrytime="00:02:35.75">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="384" swimtime="00:01:28.67" resultid="18106" heatid="19862" lane="5" entrytime="00:01:19.53" />
                <RESULT eventid="3590" points="445" swimtime="00:00:31.08" resultid="18107" heatid="19936" lane="8" entrytime="00:00:29.48" />
                <RESULT eventid="3555" points="343" reactiontime="+75" swimtime="00:01:20.08" resultid="18108" heatid="19973" lane="3" entrytime="00:01:11.81" />
                <RESULT eventid="3598" points="366" swimtime="00:01:21.25" resultid="18109" heatid="20011" lane="4" entrytime="00:01:11.33" />
                <RESULT eventid="3617" points="349" swimtime="00:00:35.58" resultid="18110" heatid="20030" lane="1" entrytime="00:00:32.04" />
                <RESULT eventid="3514" points="445" swimtime="00:00:39.03" resultid="18111" heatid="20074" lane="6" entrytime="00:00:37.97" />
                <RESULT eventid="3523" points="446" reactiontime="+77" swimtime="00:01:08.13" resultid="18112" heatid="20098" lane="4" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-09-16" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="29702" swrid="4641444" athleteid="18130">
              <RESULTS>
                <RESULT eventid="3551" points="358" swimtime="00:00:33.85" resultid="18131" heatid="19850" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="3628" points="309" reactiontime="+71" swimtime="00:01:26.62" resultid="18132" heatid="19868" lane="1" entrytime="00:01:26.40" />
                <RESULT eventid="3594" points="407" swimtime="00:00:28.20" resultid="18133" heatid="19956" lane="8" entrytime="00:00:27.48" />
                <RESULT eventid="3562" points="265" reactiontime="+76" swimtime="00:01:17.49" resultid="18134" heatid="19978" lane="2" entrytime="00:01:13.77" />
                <RESULT eventid="3605" points="330" swimtime="00:01:15.12" resultid="18135" heatid="20019" lane="3" entrytime="00:01:12.40" />
                <RESULT eventid="3613" points="371" swimtime="00:00:31.19" resultid="18136" heatid="20037" lane="2" entrytime="00:00:30.20" />
                <RESULT eventid="3519" points="328" swimtime="00:00:38.66" resultid="18137" heatid="20083" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="3530" points="360" reactiontime="+49" swimtime="00:01:05.93" resultid="18138" heatid="20108" lane="5" entrytime="00:01:01.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-10-28" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4894107" athleteid="18309">
              <RESULTS>
                <RESULT eventid="9711" points="180" reactiontime="+76" swimtime="00:03:21.61" resultid="18310" heatid="19824" lane="7" entrytime="00:03:20.09">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="170" swimtime="00:00:43.39" resultid="18311" heatid="19847" lane="8" entrytime="00:00:43.60" />
                <RESULT eventid="3594" points="199" swimtime="00:00:35.79" resultid="18312" heatid="19948" lane="7" entrytime="00:00:36.42" />
                <RESULT eventid="3512" points="155" swimtime="00:03:28.15" resultid="18313" heatid="19995" lane="8" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="152" swimtime="00:01:37.32" resultid="18314" heatid="20014" lane="6" entrytime="00:01:30.72" />
                <RESULT eventid="3613" points="94" swimtime="00:00:49.24" resultid="18315" heatid="20033" lane="6" entrytime="00:00:47.07" />
                <RESULT eventid="3519" points="134" swimtime="00:00:52.08" resultid="18316" heatid="20078" lane="7" entrytime="00:00:51.57" />
                <RESULT eventid="3530" points="168" swimtime="00:01:25.01" resultid="18317" heatid="20101" lane="3" entrytime="00:01:20.76" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-04-21" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4833278" athleteid="18139">
              <RESULTS>
                <RESULT eventid="9711" points="305" reactiontime="+61" swimtime="00:02:49.27" resultid="18140" heatid="19827" lane="1" entrytime="00:02:53.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="320" reactiontime="+63" swimtime="00:02:29.00" resultid="18141" heatid="19893" lane="6" entrytime="00:02:33.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="312" reactiontime="+71" swimtime="00:03:07.69" resultid="18142" heatid="19913" lane="6" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="294" swimtime="00:00:31.43" resultid="18143" heatid="19952" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="3605" points="261" swimtime="00:01:21.20" resultid="18144" heatid="20017" lane="1" entrytime="00:01:21.00" />
                <RESULT eventid="3613" points="243" swimtime="00:00:35.90" resultid="18145" heatid="20034" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="3519" points="312" swimtime="00:00:39.29" resultid="18146" heatid="20081" lane="2" entrytime="00:00:39.40" />
                <RESULT eventid="3530" points="325" reactiontime="+59" swimtime="00:01:08.16" resultid="18147" heatid="20106" lane="2" entrytime="00:01:07.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-04-09" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="29699" swrid="4705725" athleteid="18279">
              <RESULTS>
                <RESULT eventid="3519" points="350" swimtime="00:00:37.83" resultid="18280" heatid="20082" lane="5" entrytime="00:00:37.69" entrycourse="LCM" />
                <RESULT eventid="9711" points="349" swimtime="00:02:41.86" resultid="18281" heatid="19828" lane="5" entrytime="00:02:37.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="431" reactiontime="+90" swimtime="00:02:14.96" resultid="18282" heatid="19896" lane="1" entrytime="00:02:13.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="425" swimtime="00:00:27.81" resultid="18283" heatid="19955" lane="1" entrytime="00:00:27.77" entrycourse="LCM" />
                <RESULT eventid="3512" points="288" swimtime="00:02:49.38" resultid="18284" heatid="19998" lane="2" entrytime="00:02:43.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="305" swimtime="00:01:17.12" resultid="18285" heatid="20019" lane="7" entrytime="00:01:14.01" entrycourse="SCM" />
                <RESULT eventid="3578" points="458" reactiontime="+78" swimtime="00:04:45.31" resultid="18286" heatid="20056" lane="5" entrytime="00:04:39.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.42" />
                    <SPLIT distance="200" swimtime="00:02:20.03" />
                    <SPLIT distance="300" swimtime="00:03:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="343" reactiontime="+83" swimtime="00:01:06.96" resultid="18287" heatid="20109" lane="8" entrytime="00:01:00.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-06-20" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="41710" swrid="4879828" athleteid="18271">
              <RESULTS>
                <RESULT eventid="3639" points="340" swimtime="00:03:00.74" resultid="18272" heatid="19814" lane="5" entrytime="00:02:59.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="472" swimtime="00:02:25.10" resultid="18273" heatid="19883" lane="5" entrytime="00:02:27.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="456" swimtime="00:00:30.83" resultid="18274" heatid="19930" lane="8" entrytime="00:00:31.69" entrycourse="SCM" />
                <RESULT eventid="3505" points="332" swimtime="00:03:00.10" resultid="18275" heatid="19988" lane="8" entrytime="00:02:56.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="317" swimtime="00:01:25.23" resultid="18276" heatid="20006" lane="5" entrytime="00:01:25.11" entrycourse="SCM" />
                <RESULT eventid="3658" points="454" reactiontime="+76" swimtime="00:05:11.06" resultid="18277" heatid="20046" lane="6" entrytime="00:05:13.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="200" swimtime="00:02:32.22" />
                    <SPLIT distance="300" swimtime="00:03:52.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="444" reactiontime="+70" swimtime="00:01:08.25" resultid="18278" heatid="20095" lane="8" entrytime="00:01:07.97" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-10-06" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="29700" swrid="4781038" athleteid="18296">
              <RESULTS>
                <RESULT eventid="3551" points="284" swimtime="00:00:36.56" resultid="18297" heatid="19848" lane="5" entrytime="00:00:37.08" />
                <RESULT eventid="3628" points="259" reactiontime="+59" swimtime="00:01:31.84" resultid="18298" heatid="19868" lane="8" entrytime="00:01:26.80" />
                <RESULT eventid="3594" points="346" swimtime="00:00:29.77" resultid="18299" heatid="19953" lane="1" entrytime="00:00:29.49" />
                <RESULT eventid="3605" points="217" swimtime="00:01:26.31" resultid="18300" heatid="20017" lane="2" entrytime="00:01:19.68" />
                <RESULT eventid="3613" points="278" swimtime="00:00:34.35" resultid="18301" heatid="20036" lane="8" entrytime="00:00:32.90" />
                <RESULT eventid="3519" points="285" swimtime="00:00:40.49" resultid="18302" heatid="20081" lane="3" entrytime="00:00:38.96" />
                <RESULT eventid="3530" points="286" reactiontime="+73" swimtime="00:01:11.15" resultid="18303" heatid="20107" lane="1" entrytime="00:01:06.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-28" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="5079305" athleteid="18304">
              <RESULTS>
                <RESULT eventid="3547" points="206" swimtime="00:00:45.79" resultid="18305" heatid="19836" lane="5" entrytime="00:00:48.99" />
                <RESULT eventid="3590" points="235" swimtime="00:00:38.41" resultid="18306" heatid="19922" lane="3" entrytime="00:00:39.83" />
                <RESULT eventid="3617" points="168" swimtime="00:00:45.39" resultid="18307" heatid="20024" lane="4" entrytime="00:00:45.95" />
                <RESULT eventid="3514" points="210" swimtime="00:00:50.06" resultid="18308" heatid="20070" lane="3" entrytime="00:00:50.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-12-18" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4987131" athleteid="18202">
              <RESULTS>
                <RESULT eventid="9711" points="170" swimtime="00:03:25.57" resultid="18203" heatid="19823" lane="4" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="211" swimtime="00:02:51.14" resultid="18204" heatid="19889" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="199" swimtime="00:00:35.77" resultid="18205" heatid="19948" lane="8" entrytime="00:00:37.08" />
                <RESULT eventid="3562" points="132" swimtime="00:01:37.83" resultid="18206" heatid="19976" lane="5" entrytime="00:01:45.00" />
                <RESULT eventid="3605" points="167" swimtime="00:01:34.19" resultid="18207" heatid="20014" lane="1" entrytime="00:01:33.29" />
                <RESULT eventid="3613" points="164" swimtime="00:00:40.94" resultid="18208" heatid="20033" lane="3" entrytime="00:00:45.80" />
                <RESULT eventid="3519" points="108" swimtime="00:00:55.91" resultid="18209" heatid="20077" lane="7" entrytime="00:00:58.36" />
                <RESULT eventid="3530" points="201" reactiontime="+57" swimtime="00:01:19.96" resultid="18210" heatid="20102" lane="1" entrytime="00:01:19.64" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-11-21" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="4894093" athleteid="18087">
              <RESULTS>
                <RESULT eventid="3639" points="454" reactiontime="+60" swimtime="00:02:44.13" resultid="18088" heatid="19819" lane="1" entrytime="00:02:42.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="476" swimtime="00:02:24.62" resultid="18089" heatid="19884" lane="5" entrytime="00:02:25.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="394" swimtime="00:03:11.09" resultid="18090" heatid="19908" lane="3" entrytime="00:03:05.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="415" swimtime="00:02:47.24" resultid="18091" heatid="19990" lane="2" entrytime="00:02:43.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="397" swimtime="00:01:19.03" resultid="18092" heatid="20009" lane="5" entrytime="00:01:17.61" entrycourse="LCM" />
                <RESULT eventid="3658" points="481" reactiontime="+65" swimtime="00:05:05.20" resultid="18093" heatid="20048" lane="6" entrytime="00:05:01.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="200" swimtime="00:02:31.10" />
                    <SPLIT distance="300" swimtime="00:03:49.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" points="291" swimtime="00:03:03.69" resultid="18094" heatid="20064" lane="8" entrytime="00:02:59.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="439" swimtime="00:01:08.46" resultid="18095" heatid="20096" lane="8" entrytime="00:01:06.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-06-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="100433" swrid="4965867" athleteid="18354">
              <RESULTS>
                <RESULT eventid="3639" points="361" reactiontime="+76" swimtime="00:02:57.08" resultid="18355" heatid="19817" lane="7" entrytime="00:02:51.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="457" swimtime="00:02:26.59" resultid="18356" heatid="19885" lane="1" entrytime="00:02:24.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="419" swimtime="00:00:31.69" resultid="18357" heatid="19929" lane="2" entrytime="00:00:32.15" entrycourse="LCM" />
                <RESULT eventid="3505" points="399" swimtime="00:02:49.47" resultid="18358" heatid="19989" lane="5" entrytime="00:02:46.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="357" swimtime="00:01:21.87" resultid="18359" heatid="20009" lane="7" entrytime="00:01:19.15" entrycourse="SCM" />
                <RESULT eventid="3658" points="440" swimtime="00:05:14.27" resultid="18360" heatid="20047" lane="4" entrytime="00:05:09.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="200" swimtime="00:02:35.01" />
                    <SPLIT distance="300" swimtime="00:03:56.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="430" reactiontime="+67" swimtime="00:01:08.98" resultid="18361" heatid="20094" lane="7" entrytime="00:01:08.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-02-02" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="4987137" athleteid="18369">
              <RESULTS>
                <RESULT eventid="3639" points="319" swimtime="00:03:04.45" resultid="18370" heatid="19813" lane="7" entrytime="00:03:05.36">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="350" swimtime="00:02:40.19" resultid="18371" heatid="19880" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="308" swimtime="00:01:22.95" resultid="18372" heatid="19970" lane="2" entrytime="00:01:27.20" />
                <RESULT eventid="3505" points="315" swimtime="00:03:03.27" resultid="18373" heatid="19985" lane="1" entrytime="00:03:12.00" />
                <RESULT eventid="3617" points="310" swimtime="00:00:37.01" resultid="18374" heatid="20027" lane="7" entrytime="00:00:37.61" />
                <RESULT eventid="3658" points="363" swimtime="00:05:35.05" resultid="18375" heatid="20043" lane="1" entrytime="00:05:56.72">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.50" />
                    <SPLIT distance="200" swimtime="00:02:46.34" />
                    <SPLIT distance="300" swimtime="00:04:12.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="223" swimtime="00:00:49.13" resultid="18376" heatid="20070" lane="8" entrytime="00:00:53.46" />
                <RESULT eventid="3523" points="321" swimtime="00:01:15.98" resultid="18377" heatid="20088" lane="3" entrytime="00:01:16.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-11-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="4894110" athleteid="18384">
              <RESULTS>
                <RESULT eventid="3639" points="262" reactiontime="+70" swimtime="00:03:17.05" resultid="18385" heatid="19813" lane="8" entrytime="00:03:05.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="277" swimtime="00:00:41.47" resultid="18386" heatid="19839" lane="1" entrytime="00:00:42.54" />
                <RESULT eventid="3590" points="375" swimtime="00:00:32.90" resultid="18387" heatid="19930" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="3598" points="258" swimtime="00:01:31.24" resultid="18388" heatid="20005" lane="2" entrytime="00:01:27.90" />
                <RESULT eventid="3617" points="153" swimtime="00:00:46.85" resultid="18389" heatid="20026" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="3523" points="334" reactiontime="+69" swimtime="00:01:15.02" resultid="18390" heatid="20091" lane="7" entrytime="00:01:13.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-10-23" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="29690" swrid="4780962" athleteid="18122">
              <RESULTS>
                <RESULT eventid="3547" points="480" swimtime="00:00:34.55" resultid="18123" heatid="19842" lane="5" entrytime="00:00:35.48" entrycourse="LCM" />
                <RESULT eventid="3570" points="532" reactiontime="+82" swimtime="00:02:19.36" resultid="18124" heatid="19885" lane="7" entrytime="00:02:24.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="468" swimtime="00:00:30.55" resultid="18125" heatid="19931" lane="3" entrytime="00:00:30.92" entrycourse="LCM" />
                <RESULT eventid="3505" points="538" swimtime="00:02:33.44" resultid="18126" heatid="19990" lane="4" entrytime="00:02:41.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="512" swimtime="00:01:12.62" resultid="18127" heatid="20010" lane="6" entrytime="00:01:14.92" entrycourse="LCM" />
                <RESULT eventid="3617" points="400" swimtime="00:00:34.00" resultid="18128" heatid="20029" lane="8" entrytime="00:00:33.84" entrycourse="LCM" />
                <RESULT eventid="3523" points="491" reactiontime="+83" swimtime="00:01:05.98" resultid="18129" heatid="20096" lane="1" entrytime="00:01:06.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-08-27" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="13474" swrid="4022966" athleteid="18378">
              <RESULTS>
                <RESULT eventid="3649" points="625" swimtime="00:01:59.27" resultid="18379" heatid="19899" lane="5" entrytime="00:01:57.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="592" swimtime="00:00:24.90" resultid="18380" heatid="19958" lane="5" entrytime="00:00:24.14" entrycourse="LCM" />
                <RESULT eventid="3605" status="DNS" swimtime="00:00:00.00" resultid="18381" heatid="20022" lane="2" entrytime="00:01:01.03" entrycourse="LCM" />
                <RESULT eventid="3530" status="DNS" swimtime="00:00:00.00" resultid="18382" heatid="20112" lane="6" entrytime="00:00:52.85" entrycourse="LCM" />
                <RESULT eventid="3578" points="499" reactiontime="+72" swimtime="00:04:37.36" resultid="18383" heatid="20058" lane="3" entrytime="00:04:17.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.91" />
                    <SPLIT distance="200" swimtime="00:02:11.55" />
                    <SPLIT distance="300" swimtime="00:03:23.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15921" points="587" swimtime="00:00:24.97" resultid="20251" heatid="20121" lane="1" late="yes" />
                <RESULT eventid="15972" points="561" swimtime="00:00:25.34" resultid="20252" heatid="20123" lane="1" late="yes" />
                <RESULT eventid="15975" points="544" swimtime="00:00:25.61" resultid="20253" heatid="20125" lane="1" late="yes" />
                <RESULT eventid="15978" points="496" swimtime="00:00:26.41" resultid="20254" heatid="20127" lane="1" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-09-25" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="29695" swrid="4733821" athleteid="18422">
              <RESULTS>
                <RESULT eventid="9711" points="469" reactiontime="+78" swimtime="00:02:26.72" resultid="18423" heatid="19829" lane="3" entrytime="00:02:30.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="547" reactiontime="+68" swimtime="00:02:04.65" resultid="18424" heatid="19897" lane="1" entrytime="00:02:10.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="511" swimtime="00:00:26.15" resultid="18425" heatid="19956" lane="7" entrytime="00:00:27.24" entrycourse="LCM" />
                <RESULT eventid="3562" points="447" reactiontime="+75" swimtime="00:01:05.15" resultid="18426" heatid="19979" lane="3" entrytime="00:01:08.44" entrycourse="LCM" />
                <RESULT eventid="3613" points="514" swimtime="00:00:28.00" resultid="18427" heatid="20037" lane="6" entrytime="00:00:30.18" entrycourse="LCM" />
                <RESULT eventid="3578" points="557" reactiontime="+77" swimtime="00:04:27.36" resultid="18428" heatid="20057" lane="8" entrytime="00:04:37.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.44" />
                    <SPLIT distance="200" swimtime="00:02:10.92" />
                    <SPLIT distance="300" swimtime="00:03:20.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3588" points="403" swimtime="00:02:30.90" resultid="18429" heatid="20066" lane="5" entrytime="00:02:43.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="571" swimtime="00:00:56.53" resultid="18430" heatid="20110" lane="2" entrytime="00:00:58.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-12" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="4894100" athleteid="18211">
              <RESULTS>
                <RESULT eventid="3639" points="264" swimtime="00:03:16.46" resultid="18212" heatid="19812" lane="3" entrytime="00:03:07.44">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="246" reactiontime="+64" swimtime="00:01:42.82" resultid="18213" heatid="19857" lane="2" entrytime="00:01:36.50" />
                <RESULT eventid="3590" points="358" swimtime="00:00:33.41" resultid="18214" heatid="19927" lane="6" entrytime="00:00:33.90" />
                <RESULT eventid="3505" points="287" swimtime="00:03:09.13" resultid="18215" heatid="19987" lane="3" entrytime="00:02:58.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="273" swimtime="00:01:29.55" resultid="18216" heatid="20006" lane="6" entrytime="00:01:25.40" />
                <RESULT eventid="3617" points="199" swimtime="00:00:42.89" resultid="18217" heatid="20025" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="3514" points="280" swimtime="00:00:45.54" resultid="18218" heatid="20072" lane="7" entrytime="00:00:44.50" />
                <RESULT eventid="3523" points="297" reactiontime="+71" swimtime="00:01:18.04" resultid="18219" heatid="20091" lane="2" entrytime="00:01:13.19" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-16" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="4894094" athleteid="18096">
              <RESULTS>
                <RESULT eventid="3639" points="255" reactiontime="+77" swimtime="00:03:18.69" resultid="18097" heatid="19812" lane="6" entrytime="00:03:09.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="357" reactiontime="+73" swimtime="00:02:39.25" resultid="18098" heatid="19881" lane="2" entrytime="00:02:39.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="346" swimtime="00:00:33.77" resultid="18099" heatid="19927" lane="3" entrytime="00:00:33.79" entrycourse="LCM" />
                <RESULT eventid="3505" points="320" swimtime="00:03:02.46" resultid="18100" heatid="19987" lane="4" entrytime="00:02:57.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="305" swimtime="00:01:26.33" resultid="18101" heatid="20007" lane="2" entrytime="00:01:24.71" entrycourse="LCM" />
                <RESULT eventid="3658" points="354" reactiontime="+74" swimtime="00:05:37.78" resultid="18102" heatid="20044" lane="6" entrytime="00:05:40.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="200" swimtime="00:02:46.38" />
                    <SPLIT distance="300" swimtime="00:04:14.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="343" reactiontime="+73" swimtime="00:01:14.34" resultid="18103" heatid="20090" lane="6" entrytime="00:01:14.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-03-20" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="41709" swrid="4879825" athleteid="18175">
              <RESULTS>
                <RESULT eventid="9711" points="220" reactiontime="+85" swimtime="00:03:08.72" resultid="18176" heatid="19824" lane="6" entrytime="00:03:18.66">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="224" reactiontime="+91" swimtime="00:02:47.85" resultid="18177" heatid="19891" lane="6" entrytime="00:02:48.38">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="250" swimtime="00:00:33.15" resultid="18178" heatid="19949" lane="8" entrytime="00:00:35.38" />
                <RESULT eventid="3512" points="192" swimtime="00:03:13.90" resultid="18179" heatid="19995" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="186" swimtime="00:01:30.83" resultid="18180" heatid="20014" lane="4" entrytime="00:01:29.92" />
                <RESULT eventid="3613" points="166" swimtime="00:00:40.80" resultid="18181" heatid="20033" lane="4" entrytime="00:00:43.52" />
                <RESULT eventid="3519" points="224" swimtime="00:00:43.85" resultid="18182" heatid="20079" lane="8" entrytime="00:00:49.19" />
                <RESULT eventid="3530" points="229" swimtime="00:01:16.61" resultid="18183" heatid="20103" lane="8" entrytime="00:01:18.14" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-08-04" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4894101" athleteid="18244">
              <RESULTS>
                <RESULT eventid="9711" points="201" swimtime="00:03:14.40" resultid="18245" heatid="19824" lane="4" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="164" swimtime="00:01:46.89" resultid="18246" heatid="19864" lane="3" entrytime="00:01:45.14" />
                <RESULT eventid="3594" points="231" swimtime="00:00:34.07" resultid="18247" heatid="19949" lane="7" entrytime="00:00:35.07" />
                <RESULT eventid="3512" points="199" swimtime="00:03:11.70" resultid="18248" heatid="19995" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3613" points="143" swimtime="00:00:42.89" resultid="18249" heatid="20033" lane="7" entrytime="00:00:47.82" />
                <RESULT eventid="3578" points="237" reactiontime="+59" swimtime="00:05:55.25" resultid="18250" heatid="20052" lane="1" entrytime="00:06:04.43">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                    <SPLIT distance="200" swimtime="00:02:55.75" />
                    <SPLIT distance="300" swimtime="00:04:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="144" swimtime="00:00:50.79" resultid="18251" heatid="20078" lane="8" entrytime="00:00:52.37" />
                <RESULT eventid="3530" points="221" swimtime="00:01:17.57" resultid="18252" heatid="20102" lane="4" entrytime="00:01:18.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-07-19" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="41713" swrid="4879824" athleteid="18148">
              <RESULTS>
                <RESULT eventid="3538" points="396" reactiontime="+67" swimtime="00:03:10.67" resultid="18149" heatid="19908" lane="2" entrytime="00:03:08.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3639" points="429" swimtime="00:02:47.23" resultid="18150" heatid="19818" lane="5" entrytime="00:02:45.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="373" reactiontime="+62" swimtime="00:01:17.85" resultid="18151" heatid="19972" lane="2" entrytime="00:01:16.69" entrycourse="SCM" />
                <RESULT eventid="3598" points="364" swimtime="00:01:21.38" resultid="18152" heatid="20008" lane="4" entrytime="00:01:20.26" entrycourse="SCM" />
                <RESULT eventid="3658" points="484" reactiontime="+67" swimtime="00:05:04.54" resultid="18153" heatid="20048" lane="8" entrytime="00:05:03.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.12" />
                    <SPLIT distance="200" swimtime="00:02:31.15" />
                    <SPLIT distance="300" swimtime="00:03:49.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="401" swimtime="00:00:40.38" resultid="18154" heatid="20074" lane="8" entrytime="00:00:39.43" entrycourse="SCM" />
                <RESULT eventid="3523" points="410" reactiontime="+68" swimtime="00:01:10.08" resultid="18155" heatid="20095" lane="4" entrytime="00:01:06.99" entrycourse="SCM" />
                <RESULT eventid="3570" points="462" swimtime="00:02:26.12" resultid="18156" heatid="19884" lane="1" entrytime="00:02:26.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-06-24" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="RUS" license="41711" swrid="4879826" athleteid="18184">
              <RESULTS>
                <RESULT eventid="3551" points="285" swimtime="00:00:36.49" resultid="18185" heatid="19849" lane="8" entrytime="00:00:36.25" />
                <RESULT eventid="3628" points="318" reactiontime="+74" swimtime="00:01:25.78" resultid="18186" heatid="19868" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="3545" points="310" reactiontime="+67" swimtime="00:03:08.03" resultid="18187" heatid="19912" lane="4" entrytime="00:03:16.44">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="330" swimtime="00:00:30.25" resultid="18188" heatid="19951" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="3605" points="248" swimtime="00:01:22.58" resultid="18189" heatid="20016" lane="5" entrytime="00:01:22.90" />
                <RESULT eventid="3613" points="279" swimtime="00:00:34.32" resultid="18190" heatid="20035" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="3519" points="357" swimtime="00:00:37.59" resultid="18191" heatid="20082" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="3530" points="309" swimtime="00:01:09.36" resultid="18192" heatid="20105" lane="5" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-09-22" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="41942" swrid="4879830" athleteid="18336">
              <RESULTS>
                <RESULT eventid="3639" points="528" reactiontime="+72" swimtime="00:02:35.99" resultid="18337" heatid="19821" lane="7" entrytime="00:02:35.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="613" reactiontime="+72" swimtime="00:02:12.95" resultid="18338" heatid="19888" lane="7" entrytime="00:02:13.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="542" swimtime="00:00:29.10" resultid="18339" heatid="19936" lane="7" entrytime="00:00:28.98" entrycourse="SCM" />
                <RESULT eventid="3505" points="468" swimtime="00:02:40.69" resultid="18340" heatid="19992" lane="2" entrytime="00:02:33.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="467" swimtime="00:01:14.87" resultid="18341" heatid="20012" lane="8" entrytime="00:01:11.01" entrycourse="LCM" />
                <RESULT eventid="3658" points="560" reactiontime="+71" swimtime="00:04:49.97" resultid="18342" heatid="20050" lane="7" entrytime="00:04:44.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.92" />
                    <SPLIT distance="200" swimtime="00:02:21.98" />
                    <SPLIT distance="300" swimtime="00:03:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="532" reactiontime="+72" swimtime="00:01:04.23" resultid="18343" heatid="20099" lane="1" entrytime="00:01:02.97" entrycourse="LCM" />
                <RESULT eventid="3636" points="475" reactiontime="+77" swimtime="00:05:45.16" resultid="18344" heatid="20115" lane="6" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.58" />
                    <SPLIT distance="200" swimtime="00:02:52.56" />
                    <SPLIT distance="300" swimtime="00:04:31.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-10-08" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="29689" swrid="4781028" athleteid="18157">
              <RESULTS>
                <RESULT eventid="9711" points="276" reactiontime="+76" swimtime="00:02:55.03" resultid="18158" heatid="19826" lane="1" entrytime="00:03:00.29">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="213" reactiontime="+76" swimtime="00:01:37.97" resultid="18159" heatid="19866" lane="6" entrytime="00:01:34.18" />
                <RESULT eventid="3594" points="336" swimtime="00:00:30.06" resultid="18160" heatid="19952" lane="2" entrytime="00:00:30.25" />
                <RESULT eventid="3562" points="260" reactiontime="+74" swimtime="00:01:18.01" resultid="18161" heatid="19978" lane="7" entrytime="00:01:16.14" />
                <RESULT eventid="3605" points="258" swimtime="00:01:21.54" resultid="18162" heatid="20018" lane="8" entrytime="00:01:18.00" />
                <RESULT eventid="3613" points="296" swimtime="00:00:33.62" resultid="18163" heatid="20036" lane="6" entrytime="00:00:31.80" />
                <RESULT eventid="3519" points="237" swimtime="00:00:43.09" resultid="18164" heatid="20080" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="3530" points="314" reactiontime="+52" swimtime="00:01:08.95" resultid="18165" heatid="20106" lane="3" entrytime="00:01:07.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="27616" swrid="4621601" athleteid="18413">
              <RESULTS>
                <RESULT eventid="3639" points="486" swimtime="00:02:40.37" resultid="18414" heatid="19819" lane="4" entrytime="00:02:39.42">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="433" swimtime="00:01:25.13" resultid="18415" heatid="19861" lane="5" entrytime="00:01:22.44" />
                <RESULT eventid="3538" points="480" reactiontime="+88" swimtime="00:02:58.87" resultid="18416" heatid="19909" lane="8" entrytime="00:03:00.03">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="341" swimtime="00:01:20.24" resultid="18417" heatid="19972" lane="5" entrytime="00:01:15.98" />
                <RESULT eventid="3617" points="428" swimtime="00:00:33.26" resultid="18418" heatid="20029" lane="4" entrytime="00:00:32.19" />
                <RESULT eventid="3658" points="495" reactiontime="+69" swimtime="00:05:02.20" resultid="18419" heatid="20048" lane="2" entrytime="00:05:01.77">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="200" swimtime="00:02:27.01" />
                    <SPLIT distance="300" swimtime="00:03:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" status="DNS" swimtime="00:00:00.00" resultid="18420" heatid="20064" lane="7" entrytime="00:02:48.00" />
                <RESULT eventid="3636" points="470" reactiontime="+83" swimtime="00:05:46.55" resultid="18421" heatid="20115" lane="2" entrytime="00:05:36.88">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.22" />
                    <SPLIT distance="200" swimtime="00:02:52.75" />
                    <SPLIT distance="300" swimtime="00:04:29.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-12-27" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="25708" swrid="4413210" athleteid="18238">
              <RESULTS>
                <RESULT eventid="3639" points="555" reactiontime="+72" swimtime="00:02:33.45" resultid="18239" heatid="19821" lane="4" entrytime="00:02:34.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="552" swimtime="00:00:28.92" resultid="18240" heatid="19936" lane="6" entrytime="00:00:28.61" entrycourse="LCM" />
                <RESULT eventid="3555" points="505" reactiontime="+80" swimtime="00:01:10.37" resultid="18241" heatid="19975" lane="7" entrytime="00:01:07.91" entrycourse="LCM" />
                <RESULT eventid="3617" points="523" swimtime="00:00:31.10" resultid="18242" heatid="20031" lane="3" entrytime="00:00:29.99" entrycourse="LCM" />
                <RESULT eventid="3523" points="570" reactiontime="+79" swimtime="00:01:02.80" resultid="18243" heatid="20099" lane="6" entrytime="00:01:02.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-12-24" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="26698" swrid="4577513" athleteid="18408">
              <RESULTS>
                <RESULT eventid="3598" points="464" swimtime="00:01:15.02" resultid="18409" heatid="20011" lane="6" entrytime="00:01:12.16" />
                <RESULT eventid="3617" points="484" swimtime="00:00:31.91" resultid="18410" heatid="20030" lane="4" entrytime="00:00:31.05" />
                <RESULT eventid="3586" status="DNS" swimtime="00:00:00.00" resultid="18411" heatid="20064" lane="3" entrytime="00:02:44.90" />
                <RESULT eventid="3514" points="503" swimtime="00:00:37.45" resultid="18412" heatid="20075" lane="8" entrytime="00:00:37.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-07-13" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="26703" swrid="4577466" athleteid="18166">
              <RESULTS>
                <RESULT eventid="9711" points="546" reactiontime="+75" swimtime="00:02:19.47" resultid="18167" heatid="19832" lane="1" entrytime="00:02:20.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="567" reactiontime="+60" swimtime="00:02:03.23" resultid="18168" heatid="19897" lane="4" entrytime="00:02:07.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="454" swimtime="00:00:27.20" resultid="18169" heatid="19955" lane="8" entrytime="00:00:27.79" entrycourse="LCM" />
                <RESULT eventid="3512" points="440" swimtime="00:02:27.10" resultid="18170" heatid="20001" lane="1" entrytime="00:02:20.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="459" swimtime="00:01:07.31" resultid="18171" heatid="20021" lane="6" entrytime="00:01:05.96" entrycourse="LCM" />
                <RESULT eventid="3578" points="589" reactiontime="+72" swimtime="00:04:22.49" resultid="18172" heatid="20058" lane="8" entrytime="00:04:26.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.31" />
                    <SPLIT distance="200" swimtime="00:02:08.26" />
                    <SPLIT distance="300" swimtime="00:03:16.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="452" swimtime="00:00:34.75" resultid="18173" heatid="20083" lane="3" entrytime="00:00:35.78" entrycourse="LCM" />
                <RESULT eventid="1081" points="506" reactiontime="+76" swimtime="00:05:05.84" resultid="18174" heatid="20118" lane="3" entrytime="00:05:13.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.89" />
                    <SPLIT distance="200" swimtime="00:02:28.57" />
                    <SPLIT distance="300" swimtime="00:03:57.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-04-15" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="24813" swrid="4393961" athleteid="18362">
              <RESULTS>
                <RESULT eventid="3551" points="771" swimtime="00:00:26.21" resultid="18363" heatid="19852" lane="4" entrytime="00:00:26.40" entrycourse="LCM" />
                <RESULT eventid="3594" points="605" swimtime="00:00:24.72" resultid="18364" heatid="19957" lane="3" entrytime="00:00:25.15" entrycourse="LCM" />
                <RESULT eventid="3562" points="697" reactiontime="+54" swimtime="00:00:56.18" resultid="18365" heatid="19982" lane="4" entrytime="00:00:57.54" entrycourse="LCM" />
                <RESULT eventid="3605" points="694" swimtime="00:00:58.66" resultid="18366" heatid="20022" lane="4" entrytime="00:00:57.92" entrycourse="LCM" />
                <RESULT eventid="3613" points="662" swimtime="00:00:25.73" resultid="18367" heatid="20039" lane="3" entrytime="00:00:25.89" entrycourse="LCM" />
                <RESULT eventid="3530" points="695" reactiontime="+64" swimtime="00:00:52.95" resultid="18368" heatid="20112" lane="7" entrytime="00:00:54.27" entrycourse="LCM" />
                <RESULT eventid="15921" points="581" swimtime="00:00:25.05" resultid="20250" heatid="20121" lane="7" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-05-24" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="29691" swrid="4705726" athleteid="18327">
              <RESULTS>
                <RESULT eventid="3639" points="372" swimtime="00:02:55.28" resultid="18328" heatid="19817" lane="5" entrytime="00:02:49.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="438" swimtime="00:02:28.71" resultid="18329" heatid="19882" lane="5" entrytime="00:02:30.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="433" swimtime="00:00:31.36" resultid="18330" heatid="19931" lane="4" entrytime="00:00:30.88" entrycourse="SCM" />
                <RESULT eventid="3505" points="336" swimtime="00:02:59.41" resultid="18331" heatid="19989" lane="2" entrytime="00:02:48.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="362" swimtime="00:01:21.54" resultid="18332" heatid="20008" lane="5" entrytime="00:01:20.45" entrycourse="LCM" />
                <RESULT eventid="3658" points="405" reactiontime="+67" swimtime="00:05:23.01" resultid="18333" heatid="20046" lane="8" entrytime="00:05:16.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="200" swimtime="00:02:39.57" />
                    <SPLIT distance="300" swimtime="00:04:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="386" reactiontime="+76" swimtime="00:01:11.49" resultid="18334" heatid="20095" lane="7" entrytime="00:01:07.72" entrycourse="SCM" />
                <RESULT eventid="3636" points="325" reactiontime="+65" swimtime="00:06:31.73" resultid="18335" heatid="20114" lane="5" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.82" />
                    <SPLIT distance="200" swimtime="00:03:18.36" />
                    <SPLIT distance="300" swimtime="00:05:08.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-06-10" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" swrid="4987132" athleteid="18229">
              <RESULTS>
                <RESULT eventid="3639" points="321" reactiontime="+80" swimtime="00:03:04.20" resultid="18230" heatid="19814" lane="7" entrytime="00:03:00.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="311" swimtime="00:01:35.09" resultid="18231" heatid="19858" lane="3" entrytime="00:01:32.52" entrycourse="SCM" />
                <RESULT eventid="3538" points="326" swimtime="00:03:23.42" resultid="18232" heatid="19907" lane="1" entrytime="00:03:22.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="346" swimtime="00:02:57.68" resultid="18233" heatid="19988" lane="3" entrytime="00:02:54.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="328" swimtime="00:01:24.25" resultid="18234" heatid="20008" lane="7" entrytime="00:01:22.02" entrycourse="SCM" />
                <RESULT eventid="3658" points="384" swimtime="00:05:28.99" resultid="18235" heatid="20045" lane="2" entrytime="00:05:29.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.95" />
                    <SPLIT distance="200" swimtime="00:02:42.77" />
                    <SPLIT distance="300" swimtime="00:04:08.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="310" swimtime="00:00:44.02" resultid="18236" heatid="20072" lane="2" entrytime="00:00:43.51" entrycourse="LCM" />
                <RESULT eventid="3523" points="321" swimtime="00:01:15.99" resultid="18237" heatid="20090" lane="4" entrytime="00:01:13.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-26" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4965816" athleteid="18193">
              <RESULTS>
                <RESULT eventid="9711" points="336" reactiontime="+52" swimtime="00:02:43.98" resultid="18194" heatid="19828" lane="7" entrytime="00:02:42.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="340" reactiontime="+53" swimtime="00:02:26.10" resultid="18195" heatid="19894" lane="8" entrytime="00:02:24.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="319" swimtime="00:03:06.28" resultid="18196" heatid="19914" lane="1" entrytime="00:03:05.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="308" swimtime="00:02:45.72" resultid="18197" heatid="19998" lane="6" entrytime="00:02:42.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="281" swimtime="00:01:19.29" resultid="18198" heatid="20018" lane="6" entrytime="00:01:15.63" entrycourse="SCM" />
                <RESULT eventid="3578" points="375" reactiontime="+55" swimtime="00:05:05.10" resultid="18199" heatid="20055" lane="6" entrytime="00:05:05.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.34" />
                    <SPLIT distance="200" swimtime="00:02:32.35" />
                    <SPLIT distance="300" swimtime="00:03:51.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="295" swimtime="00:00:40.04" resultid="18200" heatid="20081" lane="7" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="3530" points="320" reactiontime="+58" swimtime="00:01:08.55" resultid="18201" heatid="20106" lane="7" entrytime="00:01:07.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="12864" points="618" reactiontime="+74" swimtime="00:03:40.94" resultid="18449" heatid="20137" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.14" />
                    <SPLIT distance="200" swimtime="00:01:50.86" />
                    <SPLIT distance="300" swimtime="00:02:47.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18378" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="18166" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="18422" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="18362" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12820" points="557" swimtime="00:04:11.85" resultid="18450" heatid="20141" lane="6" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.88" />
                    <SPLIT distance="200" swimtime="00:02:15.13" />
                    <SPLIT distance="300" swimtime="00:03:15.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18362" number="1" />
                    <RELAYPOSITION athleteid="18166" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="18378" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="18422" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="12864" points="330" reactiontime="+87" swimtime="00:04:32.34" resultid="18451" heatid="20136" lane="4" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="200" swimtime="00:02:21.24" />
                    <SPLIT distance="300" swimtime="00:03:29.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18279" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="18431" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="18193" number="3" />
                    <RELAYPOSITION athleteid="18130" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="12862" points="631" reactiontime="+60" swimtime="00:04:06.72" resultid="18452" heatid="20135" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.61" />
                    <SPLIT distance="200" swimtime="00:02:03.17" />
                    <SPLIT distance="300" swimtime="00:03:05.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18391" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="18400" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="18238" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="18336" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="3574" points="611" swimtime="00:04:33.50" resultid="18453" heatid="20139" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                    <SPLIT distance="200" swimtime="00:02:27.68" />
                    <SPLIT distance="300" swimtime="00:03:31.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18262" number="1" />
                    <RELAYPOSITION athleteid="18400" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="18391" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="18238" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="12862" points="552" reactiontime="+82" swimtime="00:04:18.00" resultid="18454" heatid="20135" lane="7" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.07" />
                    <SPLIT distance="200" swimtime="00:02:10.69" />
                    <SPLIT distance="300" swimtime="00:03:15.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18122" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="18262" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="18408" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="18345" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="3574" points="502" swimtime="00:04:52.03" resultid="18455" heatid="20138" lane="4" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.57" />
                    <SPLIT distance="200" swimtime="00:02:35.11" />
                    <SPLIT distance="300" swimtime="00:03:46.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18336" number="1" />
                    <RELAYPOSITION athleteid="18288" number="2" />
                    <RELAYPOSITION athleteid="18318" number="3" />
                    <RELAYPOSITION athleteid="18345" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="12862" points="482" reactiontime="+54" swimtime="00:04:29.99" resultid="18456" heatid="20134" lane="3" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.79" />
                    <SPLIT distance="200" swimtime="00:02:13.36" />
                    <SPLIT distance="300" swimtime="00:03:20.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18288" number="1" reactiontime="+54" />
                    <RELAYPOSITION athleteid="18271" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="18413" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="18148" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="3574" points="461" swimtime="00:05:00.54" resultid="18457" heatid="20138" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="200" swimtime="00:02:34.49" />
                    <SPLIT distance="300" swimtime="00:03:52.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18122" number="1" />
                    <RELAYPOSITION athleteid="18413" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="18148" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="18087" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SÖLL" nation="AUT" region="TLSV" clubid="14982" swrid="67828" name="Breedy Badger">
          <CONTACT city="Kufstein" email="k.leitner@kufnet.at" name="Breedy Badger" phone="05372/66157" state="AUT" street="Dr.-Karl-Erlacher-Str. 11" zip="6330" />
          <ATHLETES>
            <ATHLETE birthdate="1999-12-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38155" swrid="4736706" athleteid="18897">
              <RESULTS>
                <RESULT eventid="3590" points="476" swimtime="00:00:30.38" resultid="18898" heatid="19928" lane="7" entrytime="00:00:32.98" entrycourse="LCM" />
                <RESULT eventid="3639" points="396" swimtime="00:02:51.77" resultid="18899" heatid="19815" lane="5" entrytime="00:02:56.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="409" reactiontime="+74" swimtime="00:01:26.82" resultid="18900" heatid="19861" lane="1" entrytime="00:01:24.73" entrycourse="SCM" />
                <RESULT eventid="3555" points="407" reactiontime="+74" swimtime="00:01:15.59" resultid="18901" heatid="19973" lane="2" entrytime="00:01:12.95" entrycourse="SCM" />
                <RESULT eventid="3617" points="438" swimtime="00:00:32.99" resultid="18902" heatid="20029" lane="2" entrytime="00:00:33.23" entrycourse="SCM" />
                <RESULT eventid="3586" points="270" reactiontime="+77" swimtime="00:03:08.46" resultid="18903" heatid="20064" lane="6" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="488" reactiontime="+72" swimtime="00:01:06.12" resultid="18904" heatid="20092" lane="2" entrytime="00:01:10.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-04-18" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="39862" swrid="4826148" athleteid="18888">
              <RESULTS>
                <RESULT eventid="3639" points="376" swimtime="00:02:54.70" resultid="18889" heatid="19812" lane="5" entrytime="00:03:07.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="420" swimtime="00:01:26.03" resultid="18890" heatid="19857" lane="4" entrytime="00:01:34.73" entrycourse="LCM" />
                <RESULT eventid="3538" points="417" swimtime="00:03:07.53" resultid="18891" heatid="19907" lane="8" entrytime="00:03:24.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="368" swimtime="00:02:54.06" resultid="18892" heatid="19985" lane="5" entrytime="00:03:09.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="355" swimtime="00:01:22.04" resultid="18893" heatid="20005" lane="7" entrytime="00:01:28.03" entrycourse="LCM" />
                <RESULT eventid="3658" points="392" swimtime="00:05:26.61" resultid="18894" heatid="20044" lane="1" entrytime="00:05:45.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="200" swimtime="00:02:40.43" />
                    <SPLIT distance="300" swimtime="00:04:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="392" reactiontime="+68" swimtime="00:01:11.14" resultid="18895" heatid="20089" lane="7" entrytime="00:01:15.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-12-18" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="36390" swrid="4639767" athleteid="18848">
              <RESULTS>
                <RESULT eventid="3639" points="531" reactiontime="+76" swimtime="00:02:35.71" resultid="18849" heatid="19821" lane="8" entrytime="00:02:36.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="511" reactiontime="+75" swimtime="00:01:20.59" resultid="18850" heatid="19863" lane="6" entrytime="00:01:17.66" entrycourse="LCM" />
                <RESULT eventid="3538" points="505" reactiontime="+77" swimtime="00:02:55.85" resultid="18851" heatid="19909" lane="6" entrytime="00:02:55.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="516" swimtime="00:00:29.57" resultid="18852" heatid="19931" lane="6" entrytime="00:00:30.95" entrycourse="LCM" />
                <RESULT eventid="3505" points="520" swimtime="00:02:35.11" resultid="18853" heatid="19990" lane="3" entrytime="00:02:42.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="543" swimtime="00:01:11.24" resultid="18854" heatid="20011" lane="7" entrytime="00:01:12.52" entrycourse="LCM" />
                <RESULT eventid="3658" points="480" swimtime="00:05:05.33" resultid="18855" heatid="20047" lane="5" entrytime="00:05:09.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.73" />
                    <SPLIT distance="200" swimtime="00:02:31.19" />
                    <SPLIT distance="300" swimtime="00:03:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="524" reactiontime="+77" swimtime="00:01:04.55" resultid="18856" heatid="20096" lane="7" entrytime="00:01:06.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-10-29" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42108" swrid="5038631" athleteid="18867">
              <RESULTS>
                <RESULT eventid="3639" points="212" swimtime="00:03:31.53" resultid="18868" heatid="19811" lane="1" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="257" swimtime="00:01:41.35" resultid="18869" heatid="19854" lane="2" entrytime="00:01:48.03" entrycourse="LCM" />
                <RESULT eventid="3505" points="182" swimtime="00:03:40.19" resultid="18870" heatid="19984" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="194" swimtime="00:01:40.26" resultid="18871" heatid="20003" lane="7" entrytime="00:01:43.29" entrycourse="LCM" />
                <RESULT eventid="3658" points="188" reactiontime="+74" swimtime="00:06:57.11" resultid="18872" heatid="20041" lane="1" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.53" />
                    <SPLIT distance="200" swimtime="00:03:21.76" />
                    <SPLIT distance="300" swimtime="00:05:10.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="226" reactiontime="+75" swimtime="00:01:25.46" resultid="18873" heatid="20086" lane="6" entrytime="00:01:28.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-28" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41256" swrid="4932708" athleteid="18883">
              <RESULTS>
                <RESULT eventid="3547" points="221" swimtime="00:00:44.73" resultid="18884" heatid="19836" lane="3" entrytime="00:00:49.62" entrycourse="LCM" />
                <RESULT eventid="3590" points="240" swimtime="00:00:38.15" resultid="18885" heatid="19921" lane="4" entrytime="00:00:40.25" entrycourse="LCM" />
                <RESULT eventid="3617" points="120" swimtime="00:00:50.78" resultid="18886" heatid="20023" lane="4" entrytime="00:00:59.77" entrycourse="LCM" />
                <RESULT eventid="3514" points="233" swimtime="00:00:48.37" resultid="18887" heatid="20069" lane="4" entrytime="00:00:53.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-03-15" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38136" swrid="4826129" athleteid="18858">
              <RESULTS>
                <RESULT eventid="3639" points="321" swimtime="00:03:04.05" resultid="18859" heatid="19813" lane="4" entrytime="00:03:03.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="323" reactiontime="+60" swimtime="00:01:33.90" resultid="18860" heatid="19856" lane="3" entrytime="00:01:38.73" entrycourse="LCM" />
                <RESULT eventid="3555" points="240" reactiontime="+75" swimtime="00:01:30.13" resultid="18861" heatid="19969" lane="6" entrytime="00:01:32.55" entrycourse="LCM" />
                <RESULT eventid="3505" points="330" swimtime="00:03:00.57" resultid="18862" heatid="19986" lane="4" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="316" swimtime="00:01:25.31" resultid="18863" heatid="20007" lane="6" entrytime="00:01:24.70" entrycourse="LCM" />
                <RESULT eventid="3658" points="320" reactiontime="+74" swimtime="00:05:49.60" resultid="18864" heatid="20043" lane="6" entrytime="00:05:53.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.06" />
                    <SPLIT distance="200" swimtime="00:02:46.95" />
                    <SPLIT distance="300" swimtime="00:04:19.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="361" reactiontime="+74" swimtime="00:01:13.12" resultid="18865" heatid="20089" lane="1" entrytime="00:01:15.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCIKB" nation="AUT" region="TLSV" clubid="14167" name="Breedy Badger" shortname="SC IKB Innsbruck">
          <CONTACT email="st.opatril@aon.at" name="Breedy Badger" />
          <ATHLETES>
            <ATHLETE birthdate="2003-12-07" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="37476" swrid="4650013" athleteid="19286">
              <RESULTS>
                <RESULT eventid="3530" points="343" reactiontime="+59" swimtime="00:01:06.99" resultid="19287" heatid="20106" lane="1" entrytime="00:01:08.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-10-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="40455" swrid="4860329" athleteid="19270">
              <RESULTS>
                <RESULT eventid="9711" points="239" reactiontime="+59" swimtime="00:03:03.65" resultid="19271" heatid="19826" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="250" reactiontime="+58" swimtime="00:01:32.91" resultid="19272" heatid="19866" lane="2" entrytime="00:01:34.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-06-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="35840" swrid="4102535" athleteid="19283">
              <RESULTS>
                <RESULT eventid="3586" points="497" reactiontime="+77" swimtime="00:02:33.75" resultid="19285" heatid="20065" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-04-14" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="22971" swrid="4183036" athleteid="19256">
              <RESULTS>
                <RESULT eventid="3594" points="253" swimtime="00:00:33.02" resultid="19257" heatid="19951" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="3613" status="DNS" swimtime="00:00:00.00" resultid="19258" heatid="20035" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-11-13" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40504" swrid="4586848" athleteid="19292">
              <RESULTS>
                <RESULT eventid="3639" points="332" swimtime="00:03:02.08" resultid="19293" heatid="19813" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="312" reactiontime="+69" swimtime="00:02:46.41" resultid="19294" heatid="19880" lane="7" entrytime="00:02:46.16">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="317" swimtime="00:03:02.99" resultid="19295" heatid="19986" lane="5" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="342" swimtime="00:01:23.06" resultid="19296" heatid="20007" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="3523" points="324" reactiontime="+65" swimtime="00:01:15.75" resultid="19297" heatid="20089" lane="6" entrytime="00:01:15.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-30" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="43906" swrid="5172650" athleteid="19268">
              <RESULTS>
                <RESULT eventid="3578" points="503" reactiontime="+56" swimtime="00:04:36.70" resultid="19269" heatid="20057" lane="2" entrytime="00:04:30.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.92" />
                    <SPLIT distance="200" swimtime="00:02:13.50" />
                    <SPLIT distance="300" swimtime="00:03:24.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-02-02" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="42253" swrid="5046044" athleteid="19304">
              <RESULTS>
                <RESULT eventid="3594" points="91" swimtime="00:00:46.46" resultid="19305" heatid="19946" lane="3" entrytime="00:00:52.00" />
                <RESULT eventid="3519" points="77" swimtime="00:01:02.46" resultid="19306" heatid="20076" lane="4" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-04-10" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41193" swrid="5046041" athleteid="19276">
              <RESULTS>
                <RESULT eventid="3551" points="108" swimtime="00:00:50.38" resultid="19277" heatid="19846" lane="7" entrytime="00:01:04.98" />
                <RESULT eventid="3594" points="176" swimtime="00:00:37.26" resultid="19278" heatid="19947" lane="8" entrytime="00:00:43.98" />
                <RESULT eventid="3613" points="110" swimtime="00:00:46.70" resultid="19279" heatid="20032" lane="3" entrytime="00:00:59.97" />
                <RESULT eventid="3519" points="181" swimtime="00:00:47.14" resultid="19280" heatid="20077" lane="3" entrytime="00:00:53.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-02-17" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41533" swrid="4959522" athleteid="19313">
              <RESULTS>
                <RESULT eventid="3639" points="382" swimtime="00:02:53.75" resultid="19314" heatid="19814" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="354" swimtime="00:02:39.62" resultid="19315" heatid="19875" lane="4" entrytime="00:03:16.51">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="373" swimtime="00:00:32.96" resultid="19316" heatid="19926" lane="2" entrytime="00:00:34.54" />
                <RESULT eventid="3555" points="347" swimtime="00:01:19.73" resultid="19317" heatid="19971" lane="8" entrytime="00:01:24.15" />
                <RESULT eventid="3598" points="345" swimtime="00:01:22.79" resultid="19318" heatid="20007" lane="7" entrytime="00:01:24.90" />
                <RESULT eventid="3523" points="385" swimtime="00:01:11.56" resultid="19319" heatid="20090" lane="5" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-03-07" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" athleteid="19300">
              <RESULTS>
                <RESULT eventid="3628" points="112" reactiontime="+89" swimtime="00:02:01.23" resultid="19301" heatid="19864" lane="7" entrytime="00:02:06.00" />
                <RESULT eventid="3594" points="162" swimtime="00:00:38.33" resultid="19302" heatid="19946" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="3530" points="131" reactiontime="+87" swimtime="00:01:32.27" resultid="19303" heatid="20100" lane="2" entrytime="00:01:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-08-14" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="35334" swrid="4112389" athleteid="19241">
              <RESULTS>
                <RESULT eventid="3590" points="583" swimtime="00:00:28.40" resultid="19242" heatid="19935" lane="6" entrytime="00:00:28.63" />
                <RESULT eventid="3505" points="637" swimtime="00:02:25.05" resultid="19243" heatid="19993" lane="5" entrytime="00:02:20.52">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15921" points="576" swimtime="00:00:28.52" resultid="20194" heatid="20120" lane="1" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-03-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42248" swrid="5015011" athleteid="19230">
              <RESULTS>
                <RESULT eventid="3547" points="169" swimtime="00:00:48.93" resultid="19231" heatid="19835" lane="5" entrytime="00:00:55.08" />
                <RESULT eventid="3590" points="170" swimtime="00:00:42.79" resultid="19232" heatid="19919" lane="6" entrytime="00:00:49.96" />
                <RESULT eventid="3617" points="75" swimtime="00:00:59.34" resultid="19233" heatid="20024" lane="8" entrytime="00:00:59.41" />
                <RESULT eventid="3514" points="133" swimtime="00:00:58.34" resultid="19234" heatid="20068" lane="3" entrytime="00:01:01.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-06-10" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41184" swrid="4925052" athleteid="19223">
              <RESULTS>
                <RESULT eventid="9711" points="234" swimtime="00:03:04.84" resultid="19224" heatid="19825" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="229" reactiontime="+58" swimtime="00:02:46.66" resultid="19225" heatid="19891" lane="7" entrytime="00:02:49.31">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="219" swimtime="00:00:34.69" resultid="19226" heatid="19948" lane="4" entrytime="00:00:35.48" />
                <RESULT eventid="3613" points="149" swimtime="00:00:42.28" resultid="19227" heatid="20034" lane="1" entrytime="00:00:42.30" />
                <RESULT eventid="3578" points="242" swimtime="00:05:52.76" resultid="19228" heatid="20052" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.99" />
                    <SPLIT distance="200" swimtime="00:02:55.67" />
                    <SPLIT distance="300" swimtime="00:04:27.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="234" reactiontime="+70" swimtime="00:01:16.03" resultid="19229" heatid="20104" lane="1" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-12-14" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="37406" swrid="4478897" athleteid="19298">
              <RESULTS>
                <RESULT eventid="3523" points="509" reactiontime="+71" swimtime="00:01:05.18" resultid="19299" heatid="20095" lane="5" entrytime="00:01:07.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-30" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41187" swrid="4925054" athleteid="19235">
              <RESULTS>
                <RESULT eventid="3639" points="159" reactiontime="+85" swimtime="00:03:52.45" resultid="19236" heatid="19809" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="156" swimtime="00:03:29.82" resultid="19237" heatid="19875" lane="8" entrytime="00:04:02.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="149" swimtime="00:00:44.73" resultid="19238" heatid="19919" lane="4" entrytime="00:00:47.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-09-20" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42249" swrid="5015007" athleteid="19251">
              <RESULTS>
                <RESULT eventid="3617" points="122" swimtime="00:00:50.51" resultid="19254" heatid="20024" lane="7" entrytime="00:00:49.98" />
                <RESULT eventid="3514" points="159" swimtime="00:00:54.96" resultid="19255" heatid="20068" lane="8" entrytime="00:01:04.81" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-07-08" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42254" swrid="5015015" athleteid="19288">
              <RESULTS>
                <RESULT eventid="3621" points="145" swimtime="00:02:02.50" resultid="19289" heatid="19853" lane="3" entrytime="00:02:05.72" />
                <RESULT eventid="3590" points="119" swimtime="00:00:48.14" resultid="19290" heatid="19921" lane="7" entrytime="00:00:42.71" />
                <RESULT eventid="3523" points="157" swimtime="00:01:36.49" resultid="19291" heatid="20086" lane="8" entrytime="00:01:39.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-24" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41194" swrid="4959521" athleteid="19219">
              <RESULTS>
                <RESULT eventid="3547" points="154" swimtime="00:00:50.46" resultid="19220" heatid="19835" lane="3" entrytime="00:00:58.97" />
                <RESULT eventid="3590" points="166" swimtime="00:00:43.13" resultid="19221" heatid="19919" lane="7" entrytime="00:00:50.31" />
                <RESULT eventid="3514" points="152" swimtime="00:00:55.77" resultid="19222" heatid="20068" lane="5" entrytime="00:00:59.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-06-25" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38080" swrid="4769881" athleteid="19244">
              <RESULTS>
                <RESULT eventid="3658" points="368" swimtime="00:05:33.50" resultid="19245" heatid="20042" lane="2" entrytime="00:06:07.81">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.47" />
                    <SPLIT distance="200" swimtime="00:02:40.65" />
                    <SPLIT distance="300" swimtime="00:04:07.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="388" reactiontime="+70" swimtime="00:01:11.36" resultid="19246" heatid="20091" lane="8" entrytime="00:01:13.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-10-02" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="32903" swrid="4102644" athleteid="19239">
              <RESULTS>
                <RESULT eventid="3530" points="677" reactiontime="+67" swimtime="00:00:53.42" resultid="19240" heatid="20112" lane="3" entrytime="00:00:51.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-12-14" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="37411" swrid="4586850" athleteid="19247">
              <RESULTS>
                <RESULT eventid="3578" points="432" reactiontime="+58" swimtime="00:04:51.07" resultid="19248" heatid="20056" lane="2" entrytime="00:04:47.88">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.83" />
                    <SPLIT distance="200" swimtime="00:02:20.67" />
                    <SPLIT distance="300" swimtime="00:03:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="530" swimtime="00:00:32.95" resultid="19249" heatid="20083" lane="5" entrytime="00:00:34.80" />
                <RESULT eventid="3530" points="445" reactiontime="+71" swimtime="00:01:01.41" resultid="19250" heatid="20109" lane="1" entrytime="00:01:00.93" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-02" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41192" swrid="4959520" athleteid="19259">
              <RESULTS>
                <RESULT eventid="3547" points="223" swimtime="00:00:44.60" resultid="19260" heatid="19837" lane="4" entrytime="00:00:45.29" />
                <RESULT eventid="3590" points="256" swimtime="00:00:37.35" resultid="19261" heatid="19921" lane="2" entrytime="00:00:42.45" />
                <RESULT eventid="3617" points="130" swimtime="00:00:49.40" resultid="19262" heatid="20024" lane="6" entrytime="00:00:48.86" />
                <RESULT eventid="3514" points="309" swimtime="00:00:44.04" resultid="19263" heatid="20071" lane="8" entrytime="00:00:46.14" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-11-12" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40454" swrid="4703542" athleteid="19264">
              <RESULTS>
                <RESULT eventid="3658" points="430" reactiontime="+72" swimtime="00:05:16.61" resultid="19265" heatid="20045" lane="4" entrytime="00:05:21.55">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.97" />
                    <SPLIT distance="200" swimtime="00:02:35.20" />
                    <SPLIT distance="300" swimtime="00:03:56.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="538" swimtime="00:00:36.63" resultid="19266" heatid="20075" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="3523" points="403" reactiontime="+61" swimtime="00:01:10.48" resultid="19267" heatid="20092" lane="7" entrytime="00:01:10.97" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-03-09" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41695" swrid="5015010" athleteid="19307">
              <RESULTS>
                <RESULT comment=" - Verlassen der Schwimmlage (Zeit: 11:21)" eventid="9711" status="DSQ" swimtime="00:03:20.11" resultid="19308" heatid="19823" lane="1" />
                <RESULT eventid="3594" points="219" swimtime="00:00:34.67" resultid="19309" heatid="19947" lane="3" entrytime="00:00:39.04" />
                <RESULT eventid="3512" points="221" swimtime="00:03:04.97" resultid="19310" heatid="19994" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="220" swimtime="00:01:26.03" resultid="19311" heatid="20013" lane="2" />
                <RESULT eventid="3530" points="200" reactiontime="+64" swimtime="00:01:20.18" resultid="19312" heatid="20100" lane="1" />
                <RESULT eventid="3628" points="204" reactiontime="+69" swimtime="00:01:39.43" resultid="19784" heatid="19866" lane="1" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-07-02" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="37269" swrid="4600854" athleteid="19281">
              <RESULTS>
                <RESULT eventid="3530" points="471" reactiontime="+64" swimtime="00:01:00.25" resultid="19282" heatid="20109" lane="7" entrytime="00:01:00.68" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BLUDENZ" nation="AUT" region="VLSV" clubid="13863" name="Breedy Badger">
          <CONTACT city="Nenzing" email="mathias_eder@hotmail.com" name="Breedy Badger" street="Muttenbühel 2" zip="6710" />
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="037043" swrid="4813306" athleteid="17443">
              <RESULTS>
                <RESULT eventid="3551" status="DNS" swimtime="00:00:00.00" resultid="17444" heatid="19849" lane="5" entrytime="00:00:34.69" />
                <RESULT eventid="3628" points="425" reactiontime="+74" swimtime="00:01:17.89" resultid="17445" heatid="19869" lane="7" entrytime="00:01:23.33" />
                <RESULT eventid="3594" points="435" swimtime="00:00:27.59" resultid="17446" heatid="19955" lane="7" entrytime="00:00:27.70" />
                <RESULT eventid="3562" points="420" reactiontime="+71" swimtime="00:01:06.52" resultid="17447" heatid="19980" lane="3" entrytime="00:01:05.01" />
                <RESULT eventid="3613" points="473" swimtime="00:00:28.77" resultid="17448" heatid="20038" lane="8" entrytime="00:00:29.65" />
                <RESULT eventid="3588" points="398" reactiontime="+58" swimtime="00:02:31.49" resultid="17449" heatid="20066" lane="3" entrytime="00:02:47.05">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="382" swimtime="00:00:36.74" resultid="17450" heatid="20081" lane="4" entrytime="00:00:38.76" />
                <RESULT eventid="3530" points="424" reactiontime="+64" swimtime="00:01:02.43" resultid="17451" heatid="20109" lane="2" entrytime="00:01:00.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="038250" swrid="4520433" athleteid="17377">
              <RESULTS>
                <RESULT eventid="9711" points="270" reactiontime="+62" swimtime="00:02:56.26" resultid="17378" heatid="19824" lane="1" entrytime="00:03:21.44">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="268" reactiontime="+68" swimtime="00:01:30.76" resultid="17379" heatid="19865" lane="8" entrytime="00:01:39.06" />
                <RESULT eventid="3594" points="320" swimtime="00:00:30.56" resultid="17380" heatid="19948" lane="3" entrytime="00:00:36.19" />
                <RESULT eventid="3613" points="277" swimtime="00:00:34.40" resultid="17381" heatid="20033" lane="5" entrytime="00:00:45.47" />
                <RESULT eventid="3519" points="288" swimtime="00:00:40.35" resultid="17382" heatid="20079" lane="2" entrytime="00:00:47.15" />
                <RESULT eventid="3530" points="299" reactiontime="+60" swimtime="00:01:10.15" resultid="17383" heatid="20103" lane="1" entrytime="00:01:17.75" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="037862" swrid="4520434" athleteid="17392">
              <RESULTS>
                <RESULT eventid="9711" points="395" reactiontime="+82" swimtime="00:02:35.32" resultid="17393" heatid="19829" lane="7" entrytime="00:02:34.78">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="415" reactiontime="+81" swimtime="00:02:16.67" resultid="17394" heatid="19897" lane="8" entrytime="00:02:10.74">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="419" swimtime="00:00:27.94" resultid="17395" heatid="19956" lane="5" entrytime="00:00:26.85" />
                <RESULT eventid="3562" points="394" reactiontime="+79" swimtime="00:01:07.94" resultid="17396" heatid="19981" lane="7" entrytime="00:01:02.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="000000" swrid="5016934" athleteid="17372">
              <RESULTS>
                <RESULT eventid="3639" points="244" reactiontime="+91" swimtime="00:03:21.74" resultid="17373" heatid="19810" lane="1" entrytime="00:03:28.63">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="209" swimtime="00:00:45.54" resultid="17374" heatid="19837" lane="5" entrytime="00:00:45.63" />
                <RESULT eventid="3621" points="321" reactiontime="+71" swimtime="00:01:34.08" resultid="17375" heatid="19857" lane="1" entrytime="00:01:37.63" />
                <RESULT eventid="3590" points="287" swimtime="00:00:35.94" resultid="17376" heatid="19923" lane="5" entrytime="00:00:37.17" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="034732" swrid="4287171" athleteid="17420">
              <RESULTS>
                <RESULT eventid="3551" points="512" swimtime="00:00:30.04" resultid="17421" heatid="19851" lane="3" entrytime="00:00:30.41" />
                <RESULT eventid="3594" points="505" swimtime="00:00:26.25" resultid="17422" heatid="19957" lane="1" entrytime="00:00:26.40" />
                <RESULT eventid="3512" points="447" swimtime="00:02:26.32" resultid="17423" heatid="20000" lane="3" entrytime="00:02:22.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="485" swimtime="00:01:06.08" resultid="17424" heatid="20021" lane="2" entrytime="00:01:06.31" />
                <RESULT eventid="3519" points="463" swimtime="00:00:34.45" resultid="17425" heatid="20080" lane="4" entrytime="00:00:41.14" />
                <RESULT eventid="3530" points="516" reactiontime="+66" swimtime="00:00:58.48" resultid="17426" heatid="20110" lane="6" entrytime="00:00:58.29" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="038422" swrid="4639738" athleteid="17427">
              <RESULTS>
                <RESULT eventid="9711" points="438" swimtime="00:02:30.10" resultid="17428" heatid="19827" lane="5" entrytime="00:02:49.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="458" swimtime="00:01:15.98" resultid="17429" heatid="19868" lane="3" entrytime="00:01:24.58" />
                <RESULT eventid="3545" points="480" reactiontime="+68" swimtime="00:02:42.57" resultid="17430" heatid="19914" lane="2" entrytime="00:03:00.61">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="350" swimtime="00:00:29.67" resultid="17431" heatid="19947" lane="5" entrytime="00:00:38.32" />
                <RESULT eventid="3613" points="349" swimtime="00:00:31.85" resultid="17432" heatid="20033" lane="2" entrytime="00:00:47.76" />
                <RESULT eventid="3519" points="467" swimtime="00:00:34.36" resultid="17433" heatid="20082" lane="1" entrytime="00:00:38.52" />
                <RESULT eventid="3530" points="398" swimtime="00:01:03.77" resultid="17434" heatid="20104" lane="3" entrytime="00:01:13.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="038419" swrid="4746972" athleteid="17384">
              <RESULTS>
                <RESULT eventid="3551" points="133" swimtime="00:00:47.02" resultid="17385" heatid="19846" lane="2" entrytime="00:00:54.36" />
                <RESULT eventid="3628" points="179" reactiontime="+86" swimtime="00:01:43.85" resultid="17386" heatid="19864" lane="2" entrytime="00:01:50.24" />
                <RESULT eventid="3594" points="170" swimtime="00:00:37.71" resultid="17387" heatid="19947" lane="7" entrytime="00:00:41.94" />
                <RESULT eventid="3605" points="123" swimtime="00:01:44.27" resultid="17388" heatid="20013" lane="6" entrytime="00:01:51.76" />
                <RESULT eventid="3578" points="168" swimtime="00:06:38.13" resultid="17389" heatid="20051" lane="2" entrytime="00:07:09.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.69" />
                    <SPLIT distance="200" swimtime="00:03:13.89" />
                    <SPLIT distance="300" swimtime="00:04:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="194" swimtime="00:00:46.06" resultid="17390" heatid="20079" lane="7" entrytime="00:00:48.59" />
                <RESULT eventid="3530" points="176" swimtime="00:01:23.68" resultid="17391" heatid="20100" lane="5" entrytime="00:01:39.62" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="034726" swrid="4287174" athleteid="17435">
              <RESULTS>
                <RESULT eventid="9711" points="534" reactiontime="+61" swimtime="00:02:20.49" resultid="17436" heatid="19831" lane="3" entrytime="00:02:21.38">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="574" reactiontime="+67" swimtime="00:01:10.48" resultid="17437" heatid="19872" lane="3" entrytime="00:01:07.68" />
                <RESULT eventid="3545" points="528" reactiontime="+75" swimtime="00:02:37.49" resultid="17438" heatid="19916" lane="5" entrytime="00:02:26.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="416" reactiontime="+74" swimtime="00:01:06.71" resultid="17439" heatid="19979" lane="2" entrytime="00:01:08.88" />
                <RESULT eventid="3613" points="464" swimtime="00:00:28.97" resultid="17440" heatid="20037" lane="4" entrytime="00:00:29.76" />
                <RESULT eventid="3519" points="616" swimtime="00:00:31.33" resultid="17441" heatid="20084" lane="5" entrytime="00:00:30.57" />
                <RESULT eventid="3530" points="476" reactiontime="+64" swimtime="00:01:00.05" resultid="17442" heatid="20110" lane="3" entrytime="00:00:57.53" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="034735" swrid="4287169" athleteid="17405">
              <RESULTS>
                <RESULT eventid="9711" points="503" reactiontime="+62" swimtime="00:02:23.27" resultid="17406" heatid="19831" lane="6" entrytime="00:02:21.46">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="534" reactiontime="+63" swimtime="00:01:12.20" resultid="17407" heatid="19872" lane="6" entrytime="00:01:08.46" />
                <RESULT eventid="3594" points="537" swimtime="00:00:25.71" resultid="17408" heatid="19959" lane="6" entrytime="00:00:25.21" />
                <RESULT eventid="3613" points="487" swimtime="00:00:28.50" resultid="17409" heatid="20038" lane="7" entrytime="00:00:28.91" />
                <RESULT eventid="3519" points="604" swimtime="00:00:31.54" resultid="17410" heatid="20084" lane="3" entrytime="00:00:30.71" />
                <RESULT eventid="3530" points="572" reactiontime="+64" swimtime="00:00:56.50" resultid="17411" heatid="20112" lane="8" entrytime="00:00:54.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="000000" swrid="5148145" athleteid="17460">
              <RESULTS>
                <RESULT eventid="3551" points="104" swimtime="00:00:50.97" resultid="17461" heatid="19846" lane="1" entrytime="00:01:05.22" />
                <RESULT eventid="3594" points="137" swimtime="00:00:40.47" resultid="17462" heatid="19946" lane="6" entrytime="00:00:52.40" />
                <RESULT eventid="3519" points="128" swimtime="00:00:52.82" resultid="17463" heatid="20077" lane="6" entrytime="00:00:57.41" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="034737" swrid="4794017" athleteid="17464" />
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="000000" swrid="5148144" athleteid="17412">
              <RESULTS>
                <RESULT eventid="9711" points="160" swimtime="00:03:29.64" resultid="17413" heatid="19823" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="137" swimtime="00:03:17.43" resultid="17414" heatid="19889" lane="4" entrytime="00:03:09.67">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="147" swimtime="00:00:39.61" resultid="17415" heatid="19947" lane="1" entrytime="00:00:42.75" />
                <RESULT eventid="3512" status="DNS" swimtime="00:00:00.00" resultid="17416" heatid="19994" lane="6" entrytime="00:03:40.00" />
                <RESULT comment=" - Start vor dem Startsignal (Zeit: 11:44)" eventid="3578" reactiontime="+60" status="DSQ" swimtime="00:06:45.37" resultid="17417" heatid="20051" lane="6" entrytime="00:06:24.97">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.15" />
                    <SPLIT distance="200" swimtime="00:03:18.46" />
                    <SPLIT distance="300" swimtime="00:05:04.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="123" swimtime="00:00:53.55" resultid="17418" heatid="20076" lane="2" entrytime="00:00:58.33" />
                <RESULT eventid="3530" points="141" swimtime="00:01:30.00" resultid="17419" heatid="20100" lane="4" entrytime="00:01:30.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="000000" swrid="5046040" athleteid="17452">
              <RESULTS>
                <RESULT eventid="9711" points="146" swimtime="00:03:36.42" resultid="17453" heatid="19823" lane="7" entrytime="00:03:55.75">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="201" swimtime="00:01:39.87" resultid="17454" heatid="19864" lane="6" entrytime="00:01:49.62" />
                <RESULT eventid="3545" points="207" swimtime="00:03:35.12" resultid="17455" heatid="19911" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="192" swimtime="00:00:36.21" resultid="17456" heatid="19947" lane="2" entrytime="00:00:40.32" />
                <RESULT eventid="3613" points="118" swimtime="00:00:45.71" resultid="17457" heatid="20033" lane="1" entrytime="00:00:49.29" />
                <RESULT eventid="3519" points="211" swimtime="00:00:44.78" resultid="17458" heatid="20078" lane="6" entrytime="00:00:51.05" />
                <RESULT eventid="3530" points="167" swimtime="00:01:25.03" resultid="17459" heatid="20100" lane="3" entrytime="00:01:40.67" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="12820" points="513" swimtime="00:04:18.80" resultid="17465" heatid="20141" lane="2" entrytime="00:04:22.78">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.30" />
                    <SPLIT distance="200" swimtime="00:02:16.05" />
                    <SPLIT distance="300" swimtime="00:03:22.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17420" number="1" />
                    <RELAYPOSITION athleteid="17435" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="17392" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="17405" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12864" points="543" reactiontime="+68" swimtime="00:03:50.62" resultid="17466" heatid="20137" lane="6" entrytime="00:03:49.69">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.66" />
                    <SPLIT distance="200" swimtime="00:01:55.71" />
                    <SPLIT distance="300" swimtime="00:02:53.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17443" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="17405" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="17435" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="17420" number="4" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WITT" nation="SUI" region="ROS" clubid="16605" swrid="65667" name="Breedy Badger">
          <CONTACT city="Wittenbach" email="gabschneider@gmx.net" name="Breedy Badger" street="Grüntalstrasse 26 b" zip="9300" />
          <ATHLETES>
            <ATHLETE birthdate="2002-02-23" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="28253" swrid="4688403" athleteid="16645">
              <RESULTS>
                <RESULT eventid="3636" points="417" reactiontime="+71" swimtime="00:06:00.45" resultid="16646" heatid="20115" lane="8" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.03" />
                    <SPLIT distance="200" swimtime="00:02:58.08" />
                    <SPLIT distance="300" swimtime="00:04:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3639" points="415" reactiontime="+74" swimtime="00:02:49.09" resultid="16647" heatid="19818" lane="1" entrytime="00:02:47.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="402" reactiontime="+77" swimtime="00:01:27.29" resultid="16648" heatid="19860" lane="6" entrytime="00:01:27.54" entrycourse="LCM" />
                <RESULT eventid="3538" points="388" reactiontime="+75" swimtime="00:03:12.05" resultid="16649" heatid="19908" lane="6" entrytime="00:03:07.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="479" reactiontime="+65" swimtime="00:05:05.46" resultid="16650" heatid="20048" lane="4" entrytime="00:04:59.26">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.08" />
                    <SPLIT distance="200" swimtime="00:02:29.57" />
                    <SPLIT distance="300" swimtime="00:03:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="425" swimtime="00:00:39.63" resultid="16651" heatid="20074" lane="7" entrytime="00:00:38.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-05-09" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="45988" swrid="4894090" athleteid="16722">
              <RESULTS>
                <RESULT eventid="3639" points="298" swimtime="00:03:08.76" resultid="16723" heatid="19812" lane="1" entrytime="00:03:13.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="310" reactiontime="+72" swimtime="00:02:46.89" resultid="16724" heatid="19880" lane="6" entrytime="00:02:45.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                  </SPLITS>
                </RESULT>
                <RESULT comment=" - Verlassen der Schwimmlage (Zeit: 16:46)" eventid="3505" status="DSQ" swimtime="00:03:14.62" resultid="16725" heatid="19984" lane="2" entrytime="00:03:19.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="263" swimtime="00:01:30.60" resultid="16726" heatid="20004" lane="8" entrytime="00:01:33.27" entrycourse="LCM" />
                <RESULT eventid="3658" points="313" swimtime="00:05:51.99" resultid="16727" heatid="20043" lane="2" entrytime="00:05:54.89">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                    <SPLIT distance="200" swimtime="00:02:52.40" />
                    <SPLIT distance="300" swimtime="00:04:23.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="317" reactiontime="+60" swimtime="00:01:16.36" resultid="16728" heatid="20088" lane="7" entrytime="00:01:18.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-06-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="26263" swrid="4500016" athleteid="16630">
              <RESULTS>
                <RESULT eventid="3586" points="401" reactiontime="+72" swimtime="00:02:45.18" resultid="16631" heatid="20064" lane="4" entrytime="00:02:43.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3639" points="532" reactiontime="+75" swimtime="00:02:35.60" resultid="16632" heatid="19820" lane="7" entrytime="00:02:38.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="616" swimtime="00:02:12.72" resultid="16633" heatid="19887" lane="4" entrytime="00:02:14.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="573" swimtime="00:00:28.57" resultid="16634" heatid="19937" lane="6" entrytime="00:00:28.54" entrycourse="LCM" />
                <RESULT eventid="3555" points="486" reactiontime="+73" swimtime="00:01:11.29" resultid="16635" heatid="19974" lane="5" entrytime="00:01:09.12" entrycourse="LCM" />
                <RESULT eventid="3617" points="552" swimtime="00:00:30.56" resultid="16636" heatid="20031" lane="6" entrytime="00:00:30.23" entrycourse="LCM" />
                <RESULT eventid="3523" points="587" reactiontime="+76" swimtime="00:01:02.16" resultid="16637" heatid="20099" lane="5" entrytime="00:01:00.86" entrycourse="LCM" />
                <RESULT eventid="20145" points="592" swimtime="00:00:28.25" resultid="20149" heatid="20148" lane="4" late="yes" />
                <RESULT eventid="15921" points="579" swimtime="00:00:28.46" resultid="20266" heatid="20120" lane="8" late="yes" />
                <RESULT eventid="15972" points="538" swimtime="00:00:29.17" resultid="20267" heatid="20122" lane="8" late="yes" />
                <RESULT eventid="15975" points="501" swimtime="00:00:29.87" resultid="20268" heatid="20124" lane="8" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-04-08" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="27742" swrid="4644206" athleteid="16714">
              <RESULTS>
                <RESULT eventid="9711" points="420" reactiontime="+68" swimtime="00:02:32.15" resultid="16715" heatid="19829" lane="1" entrytime="00:02:34.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="364" reactiontime="+69" swimtime="00:01:22.00" resultid="16716" heatid="19868" lane="4" entrytime="00:01:24.10" entrycourse="LCM" />
                <RESULT eventid="3545" points="401" reactiontime="+60" swimtime="00:02:52.50" resultid="16717" heatid="19915" lane="1" entrytime="00:02:52.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="296" reactiontime="+78" swimtime="00:01:14.75" resultid="16718" heatid="19978" lane="6" entrytime="00:01:13.60" entrycourse="LCM" />
                <RESULT eventid="3605" points="331" swimtime="00:01:15.05" resultid="16719" heatid="20018" lane="7" entrytime="00:01:17.69" entrycourse="LCM" />
                <RESULT eventid="3578" points="434" reactiontime="+71" swimtime="00:04:50.56" resultid="16720" heatid="20056" lane="8" entrytime="00:04:52.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.43" />
                    <SPLIT distance="200" swimtime="00:02:22.26" />
                    <SPLIT distance="300" swimtime="00:03:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="431" reactiontime="+72" swimtime="00:05:22.76" resultid="16721" heatid="20118" lane="7" entrytime="00:05:21.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.72" />
                    <SPLIT distance="200" swimtime="00:02:38.68" />
                    <SPLIT distance="300" swimtime="00:04:10.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-11-09" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="27049" swrid="4583256" athleteid="16745">
              <RESULTS>
                <RESULT eventid="3570" points="355" swimtime="00:02:39.52" resultid="16746" heatid="19880" lane="2" entrytime="00:02:45.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="296" swimtime="00:01:24.05" resultid="16747" heatid="19970" lane="4" entrytime="00:01:24.69" entrycourse="LCM" />
                <RESULT eventid="3505" points="307" swimtime="00:03:04.92" resultid="16748" heatid="19986" lane="8" entrytime="00:03:07.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3617" points="268" swimtime="00:00:38.88" resultid="16749" heatid="20027" lane="8" entrytime="00:00:38.51" entrycourse="LCM" />
                <RESULT eventid="3586" points="328" swimtime="00:02:56.60" resultid="16750" heatid="20063" lane="3" entrytime="00:03:00.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="297" swimtime="00:01:18.03" resultid="16751" heatid="20088" lane="4" entrytime="00:01:16.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-05-09" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="27046" swrid="4583253" athleteid="16660">
              <RESULTS>
                <RESULT eventid="9711" points="420" reactiontime="+87" swimtime="00:02:32.21" resultid="16661" heatid="19828" lane="2" entrytime="00:02:39.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="450" reactiontime="+82" swimtime="00:02:13.04" resultid="16662" heatid="19895" lane="7" entrytime="00:02:16.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="410" reactiontime="+85" swimtime="00:01:07.04" resultid="16663" heatid="19979" lane="6" entrytime="00:01:08.72" />
                <RESULT eventid="3512" points="370" swimtime="00:02:35.78" resultid="16664" heatid="19999" lane="8" entrytime="00:02:35.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="369" swimtime="00:01:12.41" resultid="16665" heatid="20019" lane="4" entrytime="00:01:11.83" />
                <RESULT eventid="3578" points="499" reactiontime="+85" swimtime="00:04:37.44" resultid="16666" heatid="20056" lane="7" entrytime="00:04:49.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="200" swimtime="00:02:15.46" />
                    <SPLIT distance="300" swimtime="00:03:26.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3588" points="422" reactiontime="+82" swimtime="00:02:28.56" resultid="16667" heatid="20067" lane="8" entrytime="00:02:36.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="385" reactiontime="+80" swimtime="00:01:04.45" resultid="16668" heatid="20108" lane="8" entrytime="00:01:03.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-12-21" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="26601" swrid="4605707" athleteid="16692">
              <RESULTS>
                <RESULT eventid="3547" points="580" swimtime="00:00:32.44" resultid="16693" heatid="19844" lane="1" entrytime="00:00:33.03" entrycourse="LCM" />
                <RESULT eventid="3570" points="544" reactiontime="+87" swimtime="00:02:18.37" resultid="16694" heatid="19886" lane="7" entrytime="00:02:20.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="489" swimtime="00:00:30.10" resultid="16695" heatid="19933" lane="6" entrytime="00:00:30.26" entrycourse="LCM" />
                <RESULT eventid="3505" points="571" swimtime="00:02:30.43" resultid="16696" heatid="19993" lane="7" entrytime="00:02:30.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="562" swimtime="00:01:10.41" resultid="16697" heatid="20012" lane="3" entrytime="00:01:09.92" entrycourse="LCM" />
                <RESULT eventid="3658" points="573" reactiontime="+82" swimtime="00:04:47.78" resultid="16698" heatid="20049" lane="4" entrytime="00:04:48.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="200" swimtime="00:02:22.68" />
                    <SPLIT distance="300" swimtime="00:03:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="530" reactiontime="+73" swimtime="00:01:04.32" resultid="16699" heatid="20095" lane="2" entrytime="00:01:07.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-06-13" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="45981" swrid="4795238" athleteid="16700">
              <RESULTS>
                <RESULT eventid="1081" points="400" reactiontime="+65" swimtime="00:05:30.70" resultid="16701" heatid="20118" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.68" />
                    <SPLIT distance="200" swimtime="00:02:39.67" />
                    <SPLIT distance="300" swimtime="00:04:16.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9711" points="399" swimtime="00:02:34.79" resultid="16702" heatid="19828" lane="3" entrytime="00:02:37.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="400" reactiontime="+70" swimtime="00:02:18.43" resultid="16703" heatid="19894" lane="1" entrytime="00:02:23.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="404" swimtime="00:02:31.35" resultid="16704" heatid="19999" lane="5" entrytime="00:02:32.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="372" swimtime="00:01:12.17" resultid="16705" heatid="20020" lane="8" entrytime="00:01:11.79" entrycourse="LCM" />
                <RESULT eventid="3578" points="445" swimtime="00:04:48.25" resultid="16706" heatid="20055" lane="5" entrytime="00:04:56.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.62" />
                    <SPLIT distance="200" swimtime="00:02:22.26" />
                    <SPLIT distance="300" swimtime="00:03:36.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-08-04" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="103231" swrid="5003012" athleteid="16678">
              <RESULTS>
                <RESULT eventid="9711" points="244" reactiontime="+72" swimtime="00:03:02.37" resultid="16679" heatid="19825" lane="6" entrytime="00:03:05.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="245" swimtime="00:01:33.52" resultid="16680" heatid="19865" lane="4" entrytime="00:01:36.14" entrycourse="LCM" />
                <RESULT eventid="3545" points="265" swimtime="00:03:18.12" resultid="16681" heatid="19912" lane="5" entrytime="00:03:24.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="197" swimtime="00:01:29.15" resultid="16682" heatid="20014" lane="5" entrytime="00:01:30.03" entrycourse="LCM" />
                <RESULT eventid="3578" points="262" reactiontime="+75" swimtime="00:05:43.57" resultid="16683" heatid="20053" lane="6" entrytime="00:05:54.61">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.22" />
                    <SPLIT distance="200" swimtime="00:02:49.84" />
                    <SPLIT distance="300" swimtime="00:04:18.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="244" reactiontime="+64" swimtime="00:01:15.02" resultid="16684" heatid="20103" lane="6" entrytime="00:01:15.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-17" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="24667" swrid="4352049" athleteid="16737">
              <RESULTS>
                <RESULT eventid="3605" points="437" swimtime="00:01:08.44" resultid="16738" heatid="20020" lane="6" entrytime="00:01:10.28" entrycourse="LCM" />
                <RESULT eventid="9711" points="490" reactiontime="+69" swimtime="00:02:24.59" resultid="16739" heatid="19831" lane="8" entrytime="00:02:27.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="481" reactiontime="+71" swimtime="00:02:10.12" resultid="16740" heatid="19896" lane="6" entrytime="00:02:12.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="437" reactiontime="+70" swimtime="00:01:05.65" resultid="16741" heatid="19980" lane="2" entrytime="00:01:06.58" entrycourse="LCM" />
                <RESULT eventid="3512" points="448" swimtime="00:02:26.20" resultid="16742" heatid="20000" lane="7" entrytime="00:02:26.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="540" reactiontime="+60" swimtime="00:04:30.18" resultid="16743" heatid="20056" lane="4" entrytime="00:04:37.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                    <SPLIT distance="200" swimtime="00:02:13.15" />
                    <SPLIT distance="300" swimtime="00:03:22.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="532" reactiontime="+69" swimtime="00:05:00.80" resultid="16744" heatid="20119" lane="8" entrytime="00:05:06.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.88" />
                    <SPLIT distance="200" swimtime="00:02:26.65" />
                    <SPLIT distance="300" swimtime="00:03:52.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-14" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="28909" swrid="4705720" athleteid="16752">
              <RESULTS>
                <RESULT eventid="3639" points="381" swimtime="00:02:53.88" resultid="16753" heatid="19817" lane="8" entrytime="00:02:52.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="430" reactiontime="+73" swimtime="00:02:29.60" resultid="16754" heatid="19883" lane="7" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="418" swimtime="00:00:31.73" resultid="16755" heatid="19928" lane="6" entrytime="00:00:32.84" entrycourse="LCM" />
                <RESULT eventid="3505" points="382" swimtime="00:02:51.95" resultid="16756" heatid="19988" lane="1" entrytime="00:02:56.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="295" swimtime="00:01:27.24" resultid="16757" heatid="20007" lane="5" entrytime="00:01:23.58" entrycourse="LCM" />
                <RESULT eventid="3658" points="446" swimtime="00:05:12.79" resultid="16758" heatid="20047" lane="8" entrytime="00:05:10.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.38" />
                    <SPLIT distance="200" swimtime="00:02:35.67" />
                    <SPLIT distance="300" swimtime="00:03:55.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="423" swimtime="00:01:09.34" resultid="16759" heatid="20092" lane="5" entrytime="00:01:10.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-12" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="28908" swrid="4723808" athleteid="16606">
              <RESULTS>
                <RESULT eventid="3639" points="511" swimtime="00:02:37.79" resultid="16607" heatid="19818" lane="4" bonus="yes" entrytime="00:02:43.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="549" reactiontime="+61" swimtime="00:02:17.95" resultid="16608" heatid="19886" lane="8" entrytime="00:02:21.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="535" swimtime="00:00:29.22" resultid="16609" heatid="19933" lane="5" entrytime="00:00:30.09" entrycourse="LCM" />
                <RESULT eventid="3505" points="468" swimtime="00:02:40.74" resultid="16610" heatid="19991" lane="1" entrytime="00:02:40.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="485" swimtime="00:01:13.94" resultid="16611" heatid="20011" lane="1" entrytime="00:01:12.74" entrycourse="LCM" />
                <RESULT eventid="3658" points="509" swimtime="00:04:59.39" resultid="16612" heatid="20048" lane="3" entrytime="00:05:01.06">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="200" swimtime="00:02:26.15" />
                    <SPLIT distance="300" swimtime="00:03:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="538" reactiontime="+64" swimtime="00:01:03.99" resultid="16613" heatid="20098" lane="2" entrytime="00:01:03.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-02-07" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="29934" swrid="4725139" athleteid="16669">
              <RESULTS>
                <RESULT eventid="9711" points="424" reactiontime="+67" swimtime="00:02:31.67" resultid="16670" heatid="19829" lane="2" entrytime="00:02:34.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="384" swimtime="00:01:20.59" resultid="16671" heatid="19869" lane="3" entrytime="00:01:21.38" entrycourse="LCM" />
                <RESULT eventid="3545" points="407" reactiontime="+67" swimtime="00:02:51.66" resultid="16672" heatid="19915" lane="2" entrytime="00:02:51.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="370" reactiontime="+84" swimtime="00:01:09.35" resultid="16673" heatid="19979" lane="8" entrytime="00:01:09.64" />
                <RESULT eventid="3613" points="363" swimtime="00:00:31.43" resultid="16674" heatid="20036" lane="1" entrytime="00:00:32.87" entrycourse="LCM" />
                <RESULT eventid="3578" points="480" reactiontime="+73" swimtime="00:04:40.88" resultid="16675" heatid="20056" lane="3" entrytime="00:04:42.64">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.10" />
                    <SPLIT distance="200" swimtime="00:02:16.83" />
                    <SPLIT distance="300" swimtime="00:03:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="400" swimtime="00:00:36.19" resultid="16676" heatid="20081" lane="5" entrytime="00:00:38.89" entrycourse="LCM" />
                <RESULT eventid="1081" points="420" swimtime="00:05:25.47" resultid="16677" heatid="20117" lane="5" entrytime="00:05:34.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.44" />
                    <SPLIT distance="200" swimtime="00:02:38.01" />
                    <SPLIT distance="300" swimtime="00:04:09.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-03-17" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="45986" swrid="4894086" athleteid="16614">
              <RESULTS>
                <RESULT eventid="9711" points="264" swimtime="00:02:57.66" resultid="16615" heatid="19826" lane="8" entrytime="00:03:02.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="280" reactiontime="+78" swimtime="00:02:35.75" resultid="16616" heatid="19893" lane="2" entrytime="00:02:34.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" status="DNS" swimtime="00:00:00.00" resultid="16617" heatid="19950" lane="4" entrytime="00:00:32.61" entrycourse="LCM" />
                <RESULT eventid="3512" points="215" swimtime="00:03:06.54" resultid="16618" heatid="19994" lane="4" entrytime="00:03:18.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="202" swimtime="00:01:28.42" resultid="16619" heatid="20015" lane="7" entrytime="00:01:28.13" entrycourse="LCM" />
                <RESULT eventid="3578" points="327" swimtime="00:05:19.43" resultid="16620" heatid="20054" lane="4" entrytime="00:05:30.61">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="200" swimtime="00:02:38.08" />
                    <SPLIT distance="300" swimtime="00:04:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="297" reactiontime="+61" swimtime="00:01:10.27" resultid="16621" heatid="20105" lane="4" entrytime="00:01:09.62" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-09-18" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="28294" swrid="4688385" athleteid="16707">
              <RESULTS>
                <RESULT eventid="1081" points="332" swimtime="00:05:51.92" resultid="16708" heatid="20117" lane="3" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="200" swimtime="00:02:51.72" />
                    <SPLIT distance="300" swimtime="00:04:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9711" points="300" reactiontime="+66" swimtime="00:02:50.20" resultid="16709" heatid="19827" lane="6" entrytime="00:02:51.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="256" reactiontime="+59" swimtime="00:01:32.18" resultid="16710" heatid="19867" lane="2" entrytime="00:01:30.27" entrycourse="LCM" />
                <RESULT eventid="3545" points="306" reactiontime="+59" swimtime="00:03:08.77" resultid="16711" heatid="19913" lane="7" entrytime="00:03:14.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="327" swimtime="00:05:19.13" resultid="16712" heatid="20054" lane="5" entrytime="00:05:31.71">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.77" />
                    <SPLIT distance="200" swimtime="00:02:38.10" />
                    <SPLIT distance="300" swimtime="00:04:01.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="275" swimtime="00:00:40.97" resultid="16713" heatid="20080" lane="3" entrytime="00:00:42.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-09-16" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="28912" swrid="4723822" athleteid="16638">
              <RESULTS>
                <RESULT eventid="9711" points="258" swimtime="00:02:59.04" resultid="16639" heatid="19826" lane="3" entrytime="00:02:59.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="268" swimtime="00:02:38.01" resultid="16640" heatid="19892" lane="3" entrytime="00:02:39.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="222" swimtime="00:03:04.73" resultid="16641" heatid="19996" lane="2" entrytime="00:03:05.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="228" swimtime="00:01:24.98" resultid="16642" heatid="20016" lane="1" entrytime="00:01:25.43" entrycourse="LCM" />
                <RESULT eventid="3578" points="276" swimtime="00:05:37.70" resultid="16643" heatid="20054" lane="8" entrytime="00:05:40.18">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="200" swimtime="00:02:46.73" />
                    <SPLIT distance="300" swimtime="00:04:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="256" swimtime="00:01:13.87" resultid="16644" heatid="20104" lane="2" entrytime="00:01:13.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-05-24" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="28264" swrid="4688208" athleteid="16622">
              <RESULTS>
                <RESULT eventid="3639" points="359" swimtime="00:02:57.42" resultid="16623" heatid="19815" lane="2" entrytime="00:02:57.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="378" swimtime="00:02:36.19" resultid="16624" heatid="19882" lane="8" entrytime="00:02:36.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="314" swimtime="00:01:22.41" resultid="16625" heatid="19971" lane="1" entrytime="00:01:23.04" entrycourse="LCM" />
                <RESULT eventid="3505" points="370" swimtime="00:02:53.83" resultid="16626" heatid="19988" lane="7" entrytime="00:02:55.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="350" swimtime="00:01:22.41" resultid="16627" heatid="20008" lane="2" entrytime="00:01:21.39" entrycourse="LCM" />
                <RESULT eventid="3658" points="386" swimtime="00:05:28.20" resultid="16628" heatid="20045" lane="3" entrytime="00:05:27.66">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                    <SPLIT distance="200" swimtime="00:02:42.50" />
                    <SPLIT distance="300" swimtime="00:04:07.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="382" swimtime="00:01:11.73" resultid="16629" heatid="20091" lane="5" entrytime="00:01:12.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-10-17" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" license="24142" swrid="4327813" athleteid="16729">
              <RESULTS>
                <RESULT eventid="9711" points="528" swimtime="00:02:21.01" resultid="16730" heatid="19831" lane="5" entrytime="00:02:21.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="546" reactiontime="+72" swimtime="00:02:04.75" resultid="16731" heatid="19898" lane="7" entrytime="00:02:06.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="471" reactiontime="+76" swimtime="00:01:03.99" resultid="16732" heatid="19979" lane="5" entrytime="00:01:08.13" entrycourse="LCM" />
                <RESULT eventid="3512" points="505" swimtime="00:02:20.46" resultid="16733" heatid="20000" lane="4" entrytime="00:02:21.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="478" swimtime="00:01:06.39" resultid="16734" heatid="20021" lane="7" entrytime="00:01:06.53" entrycourse="LCM" />
                <RESULT eventid="3578" points="600" reactiontime="+77" swimtime="00:04:20.91" resultid="16735" heatid="20058" lane="7" entrytime="00:04:23.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.67" />
                    <SPLIT distance="200" swimtime="00:02:09.84" />
                    <SPLIT distance="300" swimtime="00:03:17.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="569" reactiontime="+84" swimtime="00:04:54.15" resultid="16736" heatid="20119" lane="7" entrytime="00:05:02.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                    <SPLIT distance="200" swimtime="00:02:22.39" />
                    <SPLIT distance="300" swimtime="00:03:49.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-02-17" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="SUI" license="27044" swrid="4583255" athleteid="16685">
              <RESULTS>
                <RESULT eventid="3639" points="352" reactiontime="+69" swimtime="00:02:58.63" resultid="16686" heatid="19815" lane="1" entrytime="00:02:59.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="362" reactiontime="+71" swimtime="00:01:30.41" resultid="16687" heatid="19860" lane="1" entrytime="00:01:28.68" entrycourse="LCM" />
                <RESULT eventid="3538" points="371" reactiontime="+71" swimtime="00:03:14.95" resultid="16688" heatid="19907" lane="4" entrytime="00:03:14.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="321" reactiontime="+70" swimtime="00:05:49.13" resultid="16689" heatid="20043" lane="4" entrytime="00:05:51.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.55" />
                    <SPLIT distance="200" swimtime="00:02:49.24" />
                    <SPLIT distance="300" swimtime="00:04:20.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="394" swimtime="00:00:40.62" resultid="16690" heatid="20073" lane="7" entrytime="00:00:42.07" entrycourse="LCM" />
                <RESULT eventid="3523" points="339" reactiontime="+73" swimtime="00:01:14.67" resultid="16691" heatid="20090" lane="2" entrytime="00:01:14.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="12864" points="437" swimtime="00:04:08.00" resultid="16760" heatid="20136" lane="5" entrytime="00:04:10.04">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.71" />
                    <SPLIT distance="200" swimtime="00:02:01.10" />
                    <SPLIT distance="300" swimtime="00:03:05.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16729" number="1" />
                    <RELAYPOSITION athleteid="16737" number="2" />
                    <RELAYPOSITION athleteid="16669" number="3" />
                    <RELAYPOSITION athleteid="16660" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12820" points="427" swimtime="00:04:35.19" resultid="16761" heatid="20140" lane="4" entrytime="00:04:40.02">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.26" />
                    <SPLIT distance="200" swimtime="00:02:25.83" />
                    <SPLIT distance="300" swimtime="00:03:32.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16729" number="1" />
                    <RELAYPOSITION athleteid="16669" number="2" />
                    <RELAYPOSITION athleteid="16737" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="16660" number="4" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="12862" points="565" reactiontime="+67" swimtime="00:04:16.06" resultid="16762" heatid="20135" lane="3" entrytime="00:04:19.61">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.50" />
                    <SPLIT distance="200" swimtime="00:02:05.22" />
                    <SPLIT distance="300" swimtime="00:03:08.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16630" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="16606" number="2" />
                    <RELAYPOSITION athleteid="16692" number="3" reactiontime="+11" />
                    <RELAYPOSITION athleteid="16645" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="3574" points="517" swimtime="00:04:49.13" resultid="16763" heatid="20139" lane="7" entrytime="00:04:50.53">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="200" swimtime="00:02:35.81" />
                    <SPLIT distance="300" swimtime="00:03:47.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16692" number="1" />
                    <RELAYPOSITION athleteid="16645" number="2" reactiontime="+13" />
                    <RELAYPOSITION athleteid="16630" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="16606" number="4" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WÖRGL" nation="AUT" region="TLSV" clubid="14281" swrid="71933" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2003-10-22" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="40123" swrid="4703556" athleteid="18905">
              <RESULTS>
                <RESULT eventid="3605" points="282" swimtime="00:01:19.20" resultid="18906" heatid="20019" lane="8" entrytime="00:01:14.84" entrycourse="LCM" />
                <RESULT eventid="3613" points="312" swimtime="00:00:33.05" resultid="18907" heatid="20036" lane="7" entrytime="00:00:32.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-09-23" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="40124" swrid="4797173" athleteid="18910">
              <RESULTS>
                <RESULT eventid="3628" points="333" reactiontime="+50" swimtime="00:01:24.51" resultid="18911" heatid="19868" lane="7" entrytime="00:01:26.06" entrycourse="LCM" />
                <RESULT eventid="3545" points="314" reactiontime="+49" swimtime="00:03:07.11" resultid="18912" heatid="19913" lane="4" entrytime="00:03:08.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="262" swimtime="00:00:32.67" resultid="18913" heatid="19951" lane="2" entrytime="00:00:31.76" entrycourse="LCM" />
                <RESULT eventid="3613" points="291" swimtime="00:00:33.81" resultid="18914" heatid="20034" lane="3" entrytime="00:00:36.14" entrycourse="SCM" />
                <RESULT eventid="3519" points="344" swimtime="00:00:38.05" resultid="18915" heatid="20081" lane="6" entrytime="00:00:38.98" entrycourse="LCM" />
                <RESULT eventid="3530" points="295" reactiontime="+48" swimtime="00:01:10.42" resultid="18916" heatid="20105" lane="2" entrytime="00:01:10.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="5126333" athleteid="18917">
              <RESULTS>
                <RESULT eventid="3547" points="94" swimtime="00:00:59.44" resultid="18918" heatid="19834" lane="4" entrytime="00:01:10.67" entrycourse="SCM" />
                <RESULT eventid="3590" points="103" swimtime="00:00:50.53" resultid="18919" heatid="19918" lane="5" entrytime="00:01:01.62" entrycourse="LCM" />
                <RESULT eventid="3617" points="45" swimtime="00:01:10.13" resultid="18920" heatid="20023" lane="3" entrytime="00:01:13.02" entrycourse="SCM" />
                <RESULT eventid="3514" points="128" swimtime="00:00:59.09" resultid="18921" heatid="20068" lane="2" entrytime="00:01:02.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-02-27" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="5082233" athleteid="18931">
              <RESULTS>
                <RESULT eventid="3547" points="99" swimtime="00:00:58.34" resultid="18932" heatid="19835" lane="7" entrytime="00:00:59.92" entrycourse="SCM" />
                <RESULT eventid="3590" points="103" swimtime="00:00:50.49" resultid="18933" heatid="19919" lane="1" entrytime="00:00:52.70" entrycourse="SCM" />
                <RESULT eventid="3617" points="94" swimtime="00:00:54.95" resultid="18934" heatid="20023" lane="5" entrytime="00:00:59.78" entrycourse="SCM" />
                <RESULT eventid="3514" points="128" swimtime="00:00:59.12" resultid="18935" heatid="20068" lane="7" entrytime="00:01:03.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-03-26" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40126" swrid="4959527" athleteid="18922">
              <RESULTS>
                <RESULT eventid="3547" points="518" swimtime="00:00:33.68" resultid="18923" heatid="19843" lane="4" entrytime="00:00:33.37" entrycourse="LCM" />
                <RESULT eventid="3570" points="407" reactiontime="+75" swimtime="00:02:32.34" resultid="18924" heatid="19882" lane="6" entrytime="00:02:32.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="452" swimtime="00:00:30.90" resultid="18925" heatid="19932" lane="1" entrytime="00:00:30.83" entrycourse="LCM" />
                <RESULT eventid="3505" points="425" swimtime="00:02:45.95" resultid="18926" heatid="19991" lane="3" entrytime="00:02:39.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BAMBERG" nation="GER" region="02" clubid="16764" swrid="71445" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="271055" swrid="4658084" athleteid="16838">
              <RESULTS>
                <RESULT eventid="3639" points="394" swimtime="00:02:52.06" resultid="16839" heatid="19817" lane="3" entrytime="00:02:49.94">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="375" swimtime="00:00:37.52" resultid="16840" heatid="19840" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="3570" points="446" reactiontime="+85" swimtime="00:02:27.87" resultid="16841" heatid="19884" lane="7" entrytime="00:02:26.59">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="468" swimtime="00:00:30.56" resultid="16842" heatid="19934" lane="6" entrytime="00:00:29.78" />
                <RESULT eventid="3555" points="391" reactiontime="+75" swimtime="00:01:16.62" resultid="16843" heatid="19972" lane="8" entrytime="00:01:17.38" />
                <RESULT eventid="3617" points="486" swimtime="00:00:31.88" resultid="16844" heatid="20031" lane="8" entrytime="00:00:31.04" />
                <RESULT eventid="3523" points="463" reactiontime="+80" swimtime="00:01:07.28" resultid="16845" heatid="20096" lane="2" entrytime="00:01:06.16" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="235048" swrid="4658083" athleteid="16871">
              <RESULTS>
                <RESULT eventid="3639" points="295" swimtime="00:03:09.49" resultid="16872" heatid="19814" lane="4" entrytime="00:02:59.22">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="394" swimtime="00:00:36.89" resultid="16873" heatid="19841" lane="3" entrytime="00:00:37.04" />
                <RESULT eventid="3590" points="352" swimtime="00:00:33.59" resultid="16874" heatid="19928" lane="1" entrytime="00:00:33.35" />
                <RESULT eventid="3505" points="391" swimtime="00:02:50.62" resultid="16875" heatid="19989" lane="3" entrytime="00:02:47.13">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="362" swimtime="00:01:21.54" resultid="16876" heatid="20009" lane="3" entrytime="00:01:17.79" />
                <RESULT eventid="3617" points="297" swimtime="00:00:37.55" resultid="16877" heatid="20027" lane="5" entrytime="00:00:36.68" />
                <RESULT eventid="3523" points="310" swimtime="00:01:16.87" resultid="16878" heatid="20089" lane="5" entrytime="00:01:15.42" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="294281" athleteid="16780">
              <RESULTS>
                <RESULT eventid="3628" points="285" swimtime="00:01:29.00" resultid="16781" heatid="19867" lane="5" entrytime="00:01:28.26" />
                <RESULT eventid="3545" points="305" swimtime="00:03:08.93" resultid="16782" heatid="19913" lane="2" entrytime="00:03:12.05">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="233" swimtime="00:03:01.72" resultid="16783" heatid="19996" lane="3" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment=" - Kein kontinuierliches Anschwimmen der Wende (Zeit: 10:01)" eventid="3605" status="DSQ" swimtime="00:01:26.11" resultid="16784" heatid="20016" lane="6" entrytime="00:01:24.59" />
                <RESULT eventid="3613" points="280" swimtime="00:00:34.27" resultid="16785" heatid="20035" lane="5" entrytime="00:00:33.38" />
                <RESULT eventid="3519" points="270" swimtime="00:00:41.26" resultid="16786" heatid="20080" lane="5" entrytime="00:00:42.06" />
                <RESULT eventid="3530" points="318" swimtime="00:01:08.72" resultid="16787" heatid="20106" lane="4" entrytime="00:01:07.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="249112" swrid="4658091" athleteid="16804">
              <RESULTS>
                <RESULT eventid="3547" points="396" swimtime="00:00:36.82" resultid="16805" heatid="19841" lane="1" entrytime="00:00:37.57" />
                <RESULT eventid="3570" points="399" reactiontime="+57" swimtime="00:02:33.36" resultid="16806" heatid="19881" lane="4" entrytime="00:02:36.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="459" swimtime="00:00:30.76" resultid="16807" heatid="19930" lane="5" entrytime="00:00:31.42" />
                <RESULT eventid="3505" points="295" swimtime="00:03:07.29" resultid="16808" heatid="19987" lane="8" entrytime="00:03:00.74">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="312" swimtime="00:01:25.64" resultid="16809" heatid="20007" lane="3" entrytime="00:01:24.61" />
                <RESULT eventid="3658" points="365" reactiontime="+72" swimtime="00:05:34.42" resultid="16810" heatid="20045" lane="6" entrytime="00:05:28.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="200" swimtime="00:02:44.37" />
                    <SPLIT distance="300" swimtime="00:04:10.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="409" reactiontime="+56" swimtime="00:01:10.12" resultid="16811" heatid="20093" lane="2" entrytime="00:01:09.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="271060" swrid="4658092" athleteid="16820">
              <RESULTS>
                <RESULT eventid="3639" points="282" reactiontime="+82" swimtime="00:03:12.23" resultid="16821" heatid="19813" lane="6" entrytime="00:03:04.76">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="301" reactiontime="+68" swimtime="00:01:36.08" resultid="16822" heatid="19859" lane="7" entrytime="00:01:30.42" />
                <RESULT eventid="3538" points="311" reactiontime="+70" swimtime="00:03:26.64" resultid="16823" heatid="19907" lane="2" entrytime="00:03:18.66">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="338" swimtime="00:00:34.06" resultid="16824" heatid="19927" lane="2" entrytime="00:00:33.95" />
                <RESULT eventid="3658" points="299" reactiontime="+66" swimtime="00:05:57.42" resultid="16825" heatid="20042" lane="4" entrytime="00:05:57.71">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="200" swimtime="00:02:55.61" />
                    <SPLIT distance="300" swimtime="00:04:27.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="323" swimtime="00:00:43.41" resultid="16826" heatid="20073" lane="1" entrytime="00:00:42.21" />
                <RESULT eventid="3523" points="305" reactiontime="+67" swimtime="00:01:17.35" resultid="16827" heatid="20090" lane="7" entrytime="00:01:14.97" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="329286" athleteid="16788">
              <RESULTS>
                <RESULT eventid="3639" points="389" reactiontime="+64" swimtime="00:02:52.68" resultid="16789" heatid="19816" lane="6" entrytime="00:02:53.32">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="431" swimtime="00:01:25.27" resultid="16790" heatid="19860" lane="4" entrytime="00:01:25.23" />
                <RESULT eventid="3570" points="395" reactiontime="+51" swimtime="00:02:33.93" resultid="16791" heatid="19881" lane="7" entrytime="00:02:39.58">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="425" swimtime="00:03:06.23" resultid="16792" heatid="19908" lane="5" entrytime="00:03:03.32">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="269" swimtime="00:01:26.79" resultid="16793" heatid="19970" lane="3" entrytime="00:01:25.24" />
                <RESULT eventid="3598" points="259" swimtime="00:01:31.07" resultid="16794" heatid="20007" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="3514" points="461" swimtime="00:00:38.57" resultid="16795" heatid="20074" lane="2" entrytime="00:00:38.57" />
                <RESULT eventid="3523" points="391" reactiontime="+57" swimtime="00:01:11.15" resultid="16796" heatid="20091" lane="3" entrytime="00:01:12.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="307923" athleteid="16854">
              <RESULTS>
                <RESULT eventid="3551" points="248" swimtime="00:00:38.26" resultid="16855" heatid="19848" lane="3" entrytime="00:00:38.31" />
                <RESULT eventid="3649" points="270" swimtime="00:02:37.77" resultid="16856" heatid="19892" lane="4" entrytime="00:02:37.77">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="244" swimtime="00:00:33.46" resultid="16857" heatid="19950" lane="3" entrytime="00:00:33.18" />
                <RESULT eventid="3512" points="248" swimtime="00:02:57.90" resultid="16858" heatid="19997" lane="4" entrytime="00:02:54.64">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="229" swimtime="00:01:24.79" resultid="16859" heatid="20017" lane="8" entrytime="00:01:22.03" />
                <RESULT eventid="3578" points="299" swimtime="00:05:28.94" resultid="16860" heatid="20054" lane="3" entrytime="00:05:33.16">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.96" />
                    <SPLIT distance="200" swimtime="00:02:41.60" />
                    <SPLIT distance="300" swimtime="00:04:06.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="245" swimtime="00:01:14.90" resultid="16861" heatid="20104" lane="4" entrytime="00:01:13.04" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="287819" athleteid="16862">
              <RESULTS>
                <RESULT eventid="3547" points="474" swimtime="00:00:34.69" resultid="16863" heatid="19842" lane="4" entrytime="00:00:35.23" />
                <RESULT eventid="3621" points="422" reactiontime="+77" swimtime="00:01:25.87" resultid="16864" heatid="19859" lane="4" entrytime="00:01:29.53" />
                <RESULT eventid="3538" points="426" reactiontime="+65" swimtime="00:03:06.18" resultid="16865" heatid="19909" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="407" swimtime="00:01:15.61" resultid="16866" heatid="19972" lane="1" entrytime="00:01:16.98" />
                <RESULT eventid="3505" points="429" swimtime="00:02:45.44" resultid="16867" heatid="19990" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="443" swimtime="00:01:16.24" resultid="16868" heatid="20009" lane="4" entrytime="00:01:17.11" />
                <RESULT eventid="3617" points="417" swimtime="00:00:33.54" resultid="16869" heatid="20029" lane="1" entrytime="00:00:33.52" />
                <RESULT eventid="3586" points="359" reactiontime="+66" swimtime="00:02:51.29" resultid="16870" heatid="20064" lane="2" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="152683" swrid="4124173" athleteid="16846">
              <RESULTS>
                <RESULT eventid="3551" points="548" swimtime="00:00:29.36" resultid="16847" heatid="19852" lane="6" entrytime="00:00:28.54" />
                <RESULT eventid="3649" points="546" reactiontime="+76" swimtime="00:02:04.79" resultid="16848" heatid="19898" lane="6" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="528" swimtime="00:00:25.86" resultid="16849" heatid="19959" lane="2" entrytime="00:00:25.69" />
                <RESULT eventid="3562" points="474" reactiontime="+77" swimtime="00:01:03.89" resultid="16850" heatid="19982" lane="8" entrytime="00:01:00.71" />
                <RESULT eventid="3605" points="504" swimtime="00:01:05.25" resultid="16851" heatid="20021" lane="4" entrytime="00:01:04.00" />
                <RESULT eventid="3613" points="525" swimtime="00:00:27.80" resultid="16852" heatid="20038" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="3530" points="565" reactiontime="+74" swimtime="00:00:56.73" resultid="16853" heatid="20111" lane="6" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="271059" swrid="4658093" athleteid="16812">
              <RESULTS>
                <RESULT eventid="3639" points="292" swimtime="00:03:10.02" resultid="16813" heatid="19813" lane="5" entrytime="00:03:03.83">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="283" reactiontime="+57" swimtime="00:02:52.07" resultid="16814" heatid="19879" lane="8" entrytime="00:02:52.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="323" reactiontime="+54" swimtime="00:03:24.15" resultid="16815" heatid="19906" lane="1" entrytime="00:03:30.02">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="337" swimtime="00:00:34.10" resultid="16816" heatid="19927" lane="8" entrytime="00:00:34.07" />
                <RESULT eventid="3617" points="275" swimtime="00:00:38.53" resultid="16817" heatid="20026" lane="5" entrytime="00:00:40.32" />
                <RESULT eventid="3514" points="408" swimtime="00:00:40.16" resultid="16818" heatid="20072" lane="6" entrytime="00:00:43.25" />
                <RESULT eventid="3523" points="301" reactiontime="+55" swimtime="00:01:17.69" resultid="16819" heatid="20089" lane="3" entrytime="00:01:15.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="342435" athleteid="16828">
              <RESULTS>
                <RESULT eventid="3639" points="354" reactiontime="+68" swimtime="00:02:58.26" resultid="16829" heatid="19815" lane="4" entrytime="00:02:56.53">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="384" swimtime="00:02:35.40" resultid="16830" heatid="19881" lane="3" entrytime="00:02:37.71">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="364" reactiontime="+57" swimtime="00:03:16.14" resultid="16831" heatid="19907" lane="3" entrytime="00:03:16.64">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="202" reactiontime="+84" swimtime="00:01:35.45" resultid="16832" heatid="19970" lane="8" entrytime="00:01:29.36" />
                <RESULT eventid="3617" points="299" swimtime="00:00:37.46" resultid="16833" heatid="20026" lane="3" entrytime="00:00:40.42" />
                <RESULT eventid="3658" points="338" reactiontime="+77" swimtime="00:05:43.06" resultid="16834" heatid="20044" lane="2" entrytime="00:05:42.69">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="200" swimtime="00:02:44.74" />
                    <SPLIT distance="300" swimtime="00:04:14.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" points="182" reactiontime="+75" swimtime="00:03:34.74" resultid="16835" heatid="20063" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="385" swimtime="00:00:40.94" resultid="16836" heatid="20073" lane="6" entrytime="00:00:41.41" />
                <RESULT eventid="3636" points="274" reactiontime="+77" swimtime="00:06:54.43" resultid="16837" heatid="20113" lane="4" entrytime="00:06:21.33">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.33" />
                    <SPLIT distance="200" swimtime="00:03:24.22" />
                    <SPLIT distance="300" swimtime="00:05:17.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="259900" swrid="4658096" athleteid="16797">
              <RESULTS>
                <RESULT eventid="3547" points="349" swimtime="00:00:38.43" resultid="16798" heatid="19842" lane="8" entrytime="00:00:36.04" />
                <RESULT eventid="3555" points="252" reactiontime="+77" swimtime="00:01:28.75" resultid="16799" heatid="19971" lane="6" entrytime="00:01:20.13" />
                <RESULT eventid="3505" points="313" swimtime="00:03:03.68" resultid="16800" heatid="19987" lane="6" entrytime="00:02:58.78">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="319" swimtime="00:01:25.06" resultid="16801" heatid="20009" lane="1" entrytime="00:01:19.29" />
                <RESULT eventid="3617" points="285" swimtime="00:00:38.08" resultid="16802" heatid="20028" lane="1" entrytime="00:00:35.57" />
                <RESULT eventid="3523" points="353" reactiontime="+77" swimtime="00:01:13.62" resultid="16803" heatid="20091" lane="6" entrytime="00:01:13.04" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KÖBO" nation="GER" region="02" clubid="16407" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="284231" swrid="4705009" athleteid="16429">
              <RESULTS>
                <RESULT eventid="3639" points="308" swimtime="00:03:06.64" resultid="16430" heatid="19816" lane="8" entrytime="00:02:56.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="287" swimtime="00:00:40.98" resultid="16431" heatid="19840" lane="6" entrytime="00:00:38.49" />
                <RESULT eventid="3621" points="363" reactiontime="+69" swimtime="00:01:30.31" resultid="16432" heatid="19860" lane="3" entrytime="00:01:27.39" />
                <RESULT eventid="3538" points="351" reactiontime="+82" swimtime="00:03:18.59" resultid="16433" heatid="19908" lane="7" entrytime="00:03:09.13">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="366" swimtime="00:00:33.16" resultid="16434" heatid="19929" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="3505" points="255" swimtime="00:03:16.74" resultid="16435" heatid="19988" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="257" swimtime="00:01:31.39" resultid="16436" heatid="20008" lane="8" entrytime="00:01:22.97" />
                <RESULT eventid="3658" points="286" reactiontime="+84" swimtime="00:06:02.68" resultid="16437" heatid="20040" lane="4" entrytime="00:06:44.43">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                    <SPLIT distance="200" swimtime="00:02:57.29" />
                    <SPLIT distance="300" swimtime="00:04:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="393" swimtime="00:00:40.68" resultid="16438" heatid="20074" lane="1" entrytime="00:00:39.30" />
                <RESULT eventid="3523" points="328" reactiontime="+86" swimtime="00:01:15.43" resultid="16439" heatid="20092" lane="1" entrytime="00:01:11.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="268083" swrid="4577401" athleteid="16408">
              <RESULTS>
                <RESULT eventid="3639" points="405" reactiontime="+82" swimtime="00:02:50.49" resultid="16409" heatid="19819" lane="8" entrytime="00:02:43.64">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="432" swimtime="00:01:25.21" resultid="16410" heatid="19861" lane="4" entrytime="00:01:22.01" />
                <RESULT eventid="3538" points="417" reactiontime="+71" swimtime="00:03:07.42" resultid="16411" heatid="19909" lane="2" entrytime="00:02:56.83">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="430" swimtime="00:00:31.42" resultid="16412" heatid="19934" lane="4" entrytime="00:00:29.70" />
                <RESULT eventid="3505" points="340" swimtime="00:02:58.73" resultid="16413" heatid="19991" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="380" reactiontime="+69" swimtime="00:05:29.94" resultid="16414" heatid="20044" lane="3" entrytime="00:05:39.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="200" swimtime="00:02:36.86" />
                    <SPLIT distance="300" swimtime="00:04:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" status="DNS" swimtime="00:00:00.00" resultid="16415" heatid="20063" lane="6" entrytime="00:03:03.99" />
                <RESULT eventid="3514" points="461" swimtime="00:00:38.56" resultid="16416" heatid="20074" lane="4" entrytime="00:00:37.29" />
                <RESULT eventid="3523" points="407" reactiontime="+79" swimtime="00:01:10.26" resultid="16417" heatid="20096" lane="3" entrytime="00:01:05.79" />
                <RESULT eventid="3636" points="392" reactiontime="+75" swimtime="00:06:07.91" resultid="16418" heatid="20114" lane="2" entrytime="00:06:00.92">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.64" />
                    <SPLIT distance="200" swimtime="00:03:01.41" />
                    <SPLIT distance="300" swimtime="00:04:41.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="267053" swrid="4822604" athleteid="16450">
              <RESULTS>
                <RESULT eventid="3639" points="321" swimtime="00:03:04.21" resultid="16451" heatid="19815" lane="8" entrytime="00:02:59.14">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="308" swimtime="00:00:40.06" resultid="16452" heatid="19840" lane="3" entrytime="00:00:38.33" />
                <RESULT eventid="3570" points="378" swimtime="00:02:36.20" resultid="16453" heatid="19881" lane="5" entrytime="00:02:37.31">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="403" swimtime="00:00:32.10" resultid="16454" heatid="19929" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="3555" points="242" reactiontime="+99" swimtime="00:01:29.95" resultid="16455" heatid="19970" lane="7" entrytime="00:01:28.80" />
                <RESULT eventid="3617" points="300" swimtime="00:00:37.43" resultid="16456" heatid="20027" lane="6" entrytime="00:00:37.39" />
                <RESULT eventid="3658" points="350" swimtime="00:05:39.19" resultid="16457" heatid="20044" lane="8" entrytime="00:05:50.37">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.48" />
                    <SPLIT distance="200" swimtime="00:02:47.30" />
                    <SPLIT distance="300" swimtime="00:04:17.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" points="205" swimtime="00:03:26.27" resultid="16458" heatid="20063" lane="2" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="355" swimtime="00:00:42.05" resultid="16459" heatid="20073" lane="2" entrytime="00:00:41.57" />
                <RESULT eventid="3636" points="310" swimtime="00:06:38.02" resultid="16460" heatid="20113" lane="6" entrytime="00:07:01.21">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.94" />
                    <SPLIT distance="200" swimtime="00:03:25.56" />
                    <SPLIT distance="300" swimtime="00:05:14.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="187800" swrid="4705012" athleteid="16440">
              <RESULTS>
                <RESULT eventid="3547" points="251" swimtime="00:00:42.87" resultid="16441" heatid="19840" lane="2" entrytime="00:00:38.63" />
                <RESULT eventid="3570" points="246" reactiontime="+77" swimtime="00:03:00.15" resultid="16442" heatid="19881" lane="8" entrytime="00:02:44.98">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="309" swimtime="00:00:35.09" resultid="16443" heatid="19928" lane="2" entrytime="00:00:32.86" />
                <RESULT eventid="3555" points="158" reactiontime="+69" swimtime="00:01:43.68" resultid="16444" heatid="19969" lane="7" entrytime="00:01:34.77" />
                <RESULT comment=" - Kein kontinuierliches Anschwimmen der Wende (Zeit: 9:41)" eventid="3598" status="DSQ" swimtime="00:01:34.96" resultid="16445" heatid="20006" lane="8" entrytime="00:01:26.58" />
                <RESULT eventid="3617" points="220" swimtime="00:00:41.49" resultid="16446" heatid="20027" lane="3" entrytime="00:00:37.18" />
                <RESULT eventid="3658" points="256" reactiontime="+73" swimtime="00:06:16.36" resultid="16447" heatid="20042" lane="6" entrytime="00:06:03.04">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.50" />
                    <SPLIT distance="200" swimtime="00:03:04.21" />
                    <SPLIT distance="300" swimtime="00:04:43.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="179" swimtime="00:00:52.78" resultid="16448" heatid="20070" lane="4" entrytime="00:00:46.42" />
                <RESULT eventid="3523" points="285" reactiontime="+68" swimtime="00:01:19.04" resultid="16449" heatid="20091" lane="1" entrytime="00:01:13.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="300525" swrid="4822606" athleteid="16422">
              <RESULTS>
                <RESULT eventid="9711" points="158" reactiontime="+95" swimtime="00:03:30.50" resultid="16423" heatid="19824" lane="8" entrytime="00:03:22.97">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="202" reactiontime="+82" swimtime="00:01:39.74" resultid="16424" heatid="19865" lane="2" entrytime="00:01:37.17" />
                <RESULT eventid="3649" points="163" reactiontime="+75" swimtime="00:03:06.59" resultid="16425" heatid="19890" lane="1" entrytime="00:02:56.79">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="189" swimtime="00:03:41.84" resultid="16426" heatid="19911" lane="4" entrytime="00:03:32.39">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="170" swimtime="00:00:37.72" resultid="16427" heatid="19948" lane="6" entrytime="00:00:36.25" />
                <RESULT eventid="3562" points="75" reactiontime="+85" swimtime="00:01:58.03" resultid="16428" heatid="19976" lane="3" entrytime="00:02:07.17" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="301532" swrid="4822607" athleteid="16482">
              <RESULTS>
                <RESULT eventid="9711" points="233" swimtime="00:03:05.17" resultid="16483" heatid="19826" lane="5" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="247" swimtime="00:00:38.30" resultid="16484" heatid="19848" lane="2" entrytime="00:00:40.08" />
                <RESULT eventid="3562" points="175" reactiontime="+89" swimtime="00:01:28.91" resultid="16485" heatid="19977" lane="8" entrytime="00:01:34.40" />
                <RESULT eventid="3512" points="215" swimtime="00:03:06.59" resultid="16486" heatid="19996" lane="7" entrytime="00:03:07.53">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="268027" swrid="4822616" athleteid="16461">
              <RESULTS>
                <RESULT eventid="9711" points="292" reactiontime="+75" swimtime="00:02:51.69" resultid="16462" heatid="19828" lane="8" entrytime="00:02:46.21">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="342" reactiontime="+77" swimtime="00:01:23.71" resultid="16463" heatid="19871" lane="7" entrytime="00:01:17.03" />
                <RESULT eventid="3649" points="282" reactiontime="+72" swimtime="00:02:35.45" resultid="16464" heatid="19889" lane="2" entrytime="00:03:30.01" />
                <RESULT eventid="3545" points="300" reactiontime="+82" swimtime="00:03:10.12" resultid="16465" heatid="19914" lane="7" entrytime="00:03:05.52">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="361" swimtime="00:00:29.36" resultid="16466" heatid="19954" lane="8" entrytime="00:00:28.20" />
                <RESULT eventid="3562" points="218" reactiontime="+47" swimtime="00:01:22.67" resultid="16467" heatid="19978" lane="1" entrytime="00:01:16.76" />
                <RESULT eventid="3605" points="266" swimtime="00:01:20.67" resultid="16468" heatid="20019" lane="2" entrytime="00:01:13.78" />
                <RESULT eventid="3578" points="248" reactiontime="+73" swimtime="00:05:50.11" resultid="16469" heatid="20052" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.28" />
                    <SPLIT distance="200" swimtime="00:02:53.62" />
                    <SPLIT distance="300" swimtime="00:04:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="380" reactiontime="+79" swimtime="00:01:04.76" resultid="16470" heatid="20108" lane="1" entrytime="00:01:03.63" />
                <RESULT eventid="1081" points="250" reactiontime="+48" swimtime="00:06:26.79" resultid="16471" heatid="20116" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="200" swimtime="00:03:12.48" />
                    <SPLIT distance="300" swimtime="00:05:02.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="305711" swrid="4906759" athleteid="16419">
              <RESULTS>
                <RESULT eventid="3628" points="222" reactiontime="+85" swimtime="00:01:36.73" resultid="16420" heatid="19867" lane="1" entrytime="00:01:31.24" />
                <RESULT eventid="3594" points="221" swimtime="00:00:34.57" resultid="16421" heatid="19950" lane="2" entrytime="00:00:33.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="301533" swrid="4973159" athleteid="16472">
              <RESULTS>
                <RESULT eventid="3639" points="183" reactiontime="+97" swimtime="00:03:41.86" resultid="16473" heatid="19810" lane="7" entrytime="00:03:25.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="206" swimtime="00:01:49.07" resultid="16474" heatid="19856" lane="8" entrytime="00:01:41.21" />
                <RESULT eventid="3570" points="205" reactiontime="+87" swimtime="00:03:11.41" resultid="16475" heatid="19877" lane="2" entrytime="00:02:57.15">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="270" swimtime="00:00:36.71" resultid="16476" heatid="19924" lane="5" entrytime="00:00:35.83" />
                <RESULT eventid="3555" points="114" swimtime="00:01:55.39" resultid="16477" heatid="19969" lane="1" entrytime="00:01:35.00" />
                <RESULT eventid="3617" points="150" swimtime="00:00:47.12" resultid="16478" heatid="20024" lane="3" entrytime="00:00:48.60" />
                <RESULT eventid="3658" points="203" reactiontime="+93" swimtime="00:06:46.51" resultid="16479" heatid="20041" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.38" />
                    <SPLIT distance="200" swimtime="00:03:15.74" />
                    <SPLIT distance="300" swimtime="00:05:04.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="207" swimtime="00:00:50.35" resultid="16480" heatid="20071" lane="7" entrytime="00:00:45.90" />
                <RESULT eventid="3523" points="201" swimtime="00:01:28.85" resultid="16481" heatid="20088" lane="8" entrytime="00:01:18.72" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="12820" points="212" swimtime="00:05:47.30" resultid="16487" heatid="20140" lane="3" entrytime="00:06:17.96">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="200" swimtime="00:02:58.27" />
                    <SPLIT distance="300" swimtime="00:04:20.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16461" number="1" />
                    <RELAYPOSITION athleteid="16419" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="16482" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="16422" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="3574" points="337" swimtime="00:05:33.61" resultid="16488" heatid="20138" lane="7" entrytime="00:05:41.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.13" />
                    <SPLIT distance="200" swimtime="00:03:02.38" />
                    <SPLIT distance="300" swimtime="00:04:22.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16440" number="1" />
                    <RELAYPOSITION athleteid="16429" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="16408" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="16450" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12862" points="379" swimtime="00:04:52.34" resultid="16489" heatid="20134" lane="4" entrytime="00:04:51.07">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.78" />
                    <SPLIT distance="200" swimtime="00:02:24.35" />
                    <SPLIT distance="300" swimtime="00:03:43.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16450" number="1" />
                    <RELAYPOSITION athleteid="16429" number="2" />
                    <RELAYPOSITION athleteid="16440" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="16408" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MUCSTW" nation="GER" region="02" clubid="14064" swrid="78212" name="Breedy Badger">
          <CONTACT email="200948@200941" name="Breedy Badger" />
          <ATHLETES>
            <ATHLETE birthdate="2003-04-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="368146" athleteid="18736">
              <RESULTS>
                <RESULT eventid="3605" points="342" swimtime="00:01:14.21" resultid="18737" heatid="20018" lane="2" entrytime="00:01:17.08" />
                <RESULT eventid="3613" points="321" swimtime="00:00:32.74" resultid="18738" heatid="20035" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="3519" points="348" swimtime="00:00:37.89" resultid="18739" heatid="20083" lane="8" entrytime="00:00:37.31" />
                <RESULT eventid="3530" points="409" reactiontime="+52" swimtime="00:01:03.19" resultid="18740" heatid="20107" lane="8" entrytime="00:01:07.00" />
                <RESULT eventid="1081" points="402" reactiontime="+50" swimtime="00:05:30.22" resultid="18741" heatid="20117" lane="4" entrytime="00:05:33.61">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="200" swimtime="00:02:40.60" />
                    <SPLIT distance="300" swimtime="00:04:16.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-04-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="318639" swrid="4973192" athleteid="18742">
              <RESULTS>
                <RESULT eventid="3578" points="545" swimtime="00:04:29.40" resultid="18743" heatid="20057" lane="5" entrytime="00:04:29.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.97" />
                    <SPLIT distance="200" swimtime="00:02:12.25" />
                    <SPLIT distance="300" swimtime="00:03:21.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3588" points="406" reactiontime="+75" swimtime="00:02:30.55" resultid="18744" heatid="20067" lane="1" entrytime="00:02:35.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="476" swimtime="00:01:00.07" resultid="18745" heatid="20109" lane="3" entrytime="00:00:59.76" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ZIRL" nation="AUT" region="TLSV" clubid="14824" swrid="68100" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2008-06-03" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43435" swrid="5101386" athleteid="18782">
              <RESULTS>
                <RESULT eventid="3590" points="150" swimtime="00:00:44.57" resultid="18783" heatid="19918" lane="4" entrytime="00:00:54.30" />
                <RESULT eventid="3514" points="172" swimtime="00:00:53.50" resultid="18784" heatid="20068" lane="6" entrytime="00:01:01.83" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-03" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42244" swrid="5015021" athleteid="18785">
              <RESULTS>
                <RESULT eventid="3547" points="367" swimtime="00:00:37.79" resultid="18786" heatid="19840" lane="5" entrytime="00:00:38.13" />
                <RESULT eventid="3590" points="347" swimtime="00:00:33.76" resultid="18787" heatid="19926" lane="5" entrytime="00:00:34.43" />
                <RESULT eventid="3617" points="262" swimtime="00:00:39.14" resultid="18788" heatid="20025" lane="7" entrytime="00:00:44.59" />
                <RESULT eventid="3514" points="331" swimtime="00:00:43.06" resultid="18789" heatid="20071" lane="1" entrytime="00:00:45.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="33649" swrid="4102529" athleteid="18790">
              <RESULTS>
                <RESULT eventid="9711" points="592" reactiontime="+70" swimtime="00:02:15.71" resultid="18791" heatid="19832" lane="2" entrytime="00:02:13.73">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="537" swimtime="00:02:17.64" resultid="18792" heatid="20001" lane="4" entrytime="00:02:13.05">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="626" reactiontime="+71" swimtime="00:04:17.24" resultid="18793" heatid="20058" lane="5" entrytime="00:04:15.13">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.15" />
                    <SPLIT distance="200" swimtime="00:02:06.13" />
                    <SPLIT distance="300" swimtime="00:03:12.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="582" reactiontime="+72" swimtime="00:04:52.00" resultid="18794" heatid="20119" lane="5" entrytime="00:04:41.98">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                    <SPLIT distance="200" swimtime="00:02:22.32" />
                    <SPLIT distance="300" swimtime="00:03:47.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-10-14" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41148" swrid="4797190" athleteid="18795">
              <RESULTS>
                <RESULT eventid="3628" points="257" swimtime="00:01:32.06" resultid="18796" heatid="19866" lane="3" entrytime="00:01:33.91" />
                <RESULT eventid="3545" points="256" swimtime="00:03:20.37" resultid="18797" heatid="19912" lane="6" entrytime="00:03:25.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="147" swimtime="00:01:34.25" resultid="18798" heatid="19977" lane="1" entrytime="00:01:33.23" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-04" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41145" swrid="4902510" athleteid="18775">
              <RESULTS>
                <RESULT eventid="3621" points="337" reactiontime="+84" swimtime="00:01:32.53" resultid="18776" heatid="19858" lane="2" entrytime="00:01:33.95" />
                <RESULT eventid="3538" points="343" reactiontime="+85" swimtime="00:03:20.09" resultid="18777" heatid="19907" lane="7" entrytime="00:03:18.85">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="325" swimtime="00:00:34.50" resultid="18778" heatid="19925" lane="8" entrytime="00:00:35.54" />
                <RESULT eventid="3617" points="259" swimtime="00:00:39.32" resultid="18779" heatid="20026" lane="7" entrytime="00:00:40.88" />
                <RESULT eventid="3514" points="333" swimtime="00:00:42.96" resultid="18780" heatid="20072" lane="1" entrytime="00:00:44.53" />
                <RESULT eventid="3523" points="271" swimtime="00:01:20.45" resultid="18781" heatid="20087" lane="2" entrytime="00:01:21.31" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LEUT" nation="AUT" region="TLSV" clubid="14941" swrid="68099" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2006-09-11" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="RUS" license="43203" swrid="5101382" athleteid="18805">
              <RESULTS>
                <RESULT eventid="3551" points="171" swimtime="00:00:43.27" resultid="18806" heatid="19846" lane="5" entrytime="00:00:46.31" entrycourse="LCM" />
                <RESULT eventid="3594" points="181" swimtime="00:00:36.91" resultid="18807" heatid="19947" lane="4" entrytime="00:00:38.01" entrycourse="LCM" />
                <RESULT eventid="3613" points="115" swimtime="00:00:46.12" resultid="18808" heatid="20032" lane="5" entrytime="00:00:51.63" entrycourse="LCM" />
                <RESULT eventid="3519" points="160" swimtime="00:00:49.10" resultid="18809" heatid="20078" lane="5" entrytime="00:00:50.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-09-29" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" athleteid="18799">
              <RESULTS>
                <RESULT eventid="3551" points="86" swimtime="00:00:54.33" resultid="19788" heatid="19845" lane="4" />
                <RESULT eventid="3594" points="98" swimtime="00:00:45.35" resultid="19789" heatid="19945" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-12" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43204" swrid="5071976" athleteid="18831">
              <RESULTS>
                <RESULT eventid="3547" points="151" swimtime="00:00:50.78" resultid="18832" heatid="19836" lane="4" entrytime="00:00:48.11" entrycourse="SCM" />
                <RESULT eventid="3590" points="227" swimtime="00:00:38.88" resultid="18833" heatid="19922" lane="6" entrytime="00:00:39.93" entrycourse="SCM" />
                <RESULT eventid="3617" points="142" swimtime="00:00:47.97" resultid="18834" heatid="20024" lane="5" entrytime="00:00:46.33" entrycourse="SCM" />
                <RESULT eventid="3514" points="124" swimtime="00:00:59.65" resultid="18835" heatid="20069" lane="7" entrytime="00:00:56.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2009-10-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43597" athleteid="18810">
              <RESULTS>
                <RESULT eventid="3547" points="34" swimtime="00:01:22.88" resultid="18811" heatid="19833" lane="7" />
                <RESULT eventid="3590" points="27" swimtime="00:01:18.20" resultid="18812" heatid="19917" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-09-11" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43200" swrid="5101383" athleteid="18813">
              <RESULTS>
                <RESULT eventid="3547" points="135" swimtime="00:00:52.62" resultid="18814" heatid="19836" lane="6" entrytime="00:00:49.97" entrycourse="SCM" />
                <RESULT eventid="3590" points="113" swimtime="00:00:49.07" resultid="18815" heatid="19920" lane="7" entrytime="00:00:45.26" entrycourse="SCM" />
                <RESULT eventid="3617" points="58" swimtime="00:01:04.73" resultid="18816" heatid="20024" lane="1" entrytime="00:00:55.68" entrycourse="SCM" />
                <RESULT eventid="3514" points="89" swimtime="00:01:06.62" resultid="18817" heatid="20069" lane="8" entrytime="00:00:57.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-06-25" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="42271" swrid="5015018" athleteid="18828">
              <RESULTS>
                <RESULT eventid="3613" points="97" swimtime="00:00:48.68" resultid="18829" heatid="20032" lane="4" entrytime="00:00:50.89" entrycourse="LCM" />
                <RESULT eventid="3519" points="116" swimtime="00:00:54.67" resultid="18830" heatid="20077" lane="1" entrytime="00:00:58.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-05-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="39689" swrid="4925059" athleteid="18818">
              <RESULTS>
                <RESULT eventid="3639" points="298" swimtime="00:03:08.86" resultid="18819" heatid="19813" lane="1" entrytime="00:03:05.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="316" swimtime="00:01:34.55" resultid="18820" heatid="19857" lane="3" entrytime="00:01:35.16" entrycourse="SCM" />
                <RESULT eventid="3570" points="307" reactiontime="+79" swimtime="00:02:47.31" resultid="18821" heatid="19880" lane="1" entrytime="00:02:47.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="299" reactiontime="+79" swimtime="00:03:29.46" resultid="18822" heatid="19905" lane="7" entrytime="00:03:50.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="268" swimtime="00:01:30.11" resultid="18823" heatid="20006" lane="7" entrytime="00:01:25.89" entrycourse="SCM" />
                <RESULT eventid="3658" points="314" reactiontime="+82" swimtime="00:05:51.52" resultid="18824" heatid="20044" lane="7" entrytime="00:05:43.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.63" />
                    <SPLIT distance="200" swimtime="00:02:52.45" />
                    <SPLIT distance="300" swimtime="00:04:25.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3636" points="263" reactiontime="+75" swimtime="00:07:00.52" resultid="18825" heatid="20113" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.50" />
                    <SPLIT distance="200" swimtime="00:03:33.80" />
                    <SPLIT distance="300" swimtime="00:05:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="306" swimtime="00:01:17.19" resultid="18826" heatid="20090" lane="8" entrytime="00:01:15.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-11-20" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="32734" swrid="4104206" athleteid="18827" />
            <ATHLETE birthdate="2006-11-05" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43195" swrid="5082238" athleteid="18802">
              <RESULTS>
                <RESULT eventid="3547" points="114" swimtime="00:00:55.75" resultid="18803" heatid="19835" lane="4" entrytime="00:00:54.96" entrycourse="SCM" />
                <RESULT eventid="3590" points="109" swimtime="00:00:49.61" resultid="18804" heatid="19919" lane="3" entrytime="00:00:48.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="12862" points="205" swimtime="00:05:59.05" resultid="18836" heatid="20134" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.29" />
                    <SPLIT distance="200" swimtime="00:02:51.60" />
                    <SPLIT distance="300" swimtime="00:04:42.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18827" number="1" />
                    <RELAYPOSITION athleteid="18831" number="2" />
                    <RELAYPOSITION athleteid="18813" number="3" />
                    <RELAYPOSITION athleteid="18818" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="BRUNECK" nation="ITA" clubid="12874" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5164030" athleteid="17085">
              <RESULTS>
                <RESULT eventid="3547" points="141" swimtime="00:00:51.92" resultid="17086" heatid="19833" lane="2" />
                <RESULT eventid="3590" points="144" swimtime="00:00:45.18" resultid="17087" heatid="19918" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4911986" athleteid="16956">
              <RESULTS>
                <RESULT eventid="3547" points="234" swimtime="00:00:43.86" resultid="16957" heatid="19839" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="3621" points="241" swimtime="00:01:43.52" resultid="16958" heatid="19855" lane="5" entrytime="00:01:42.00" />
                <RESULT eventid="3538" points="232" reactiontime="+75" swimtime="00:03:48.01" resultid="16959" heatid="19906" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="272" swimtime="00:00:36.58" resultid="16960" heatid="19924" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" athleteid="19785">
              <RESULTS>
                <RESULT eventid="3547" points="133" swimtime="00:00:52.94" resultid="19786" heatid="19834" lane="1" />
                <RESULT eventid="3590" points="140" swimtime="00:00:45.63" resultid="19787" heatid="19918" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5093619" athleteid="16974">
              <RESULTS>
                <RESULT eventid="3547" points="155" swimtime="00:00:50.30" resultid="16975" heatid="19838" lane="3" entrytime="00:00:44.00" />
                <RESULT eventid="3570" points="182" swimtime="00:03:19.36" resultid="16976" heatid="19875" lane="5" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="207" swimtime="00:00:40.07" resultid="16977" heatid="19922" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4994491" athleteid="16936">
              <RESULTS>
                <RESULT eventid="3551" points="142" swimtime="00:00:46.05" resultid="16937" heatid="19846" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="3649" points="228" reactiontime="+89" swimtime="00:02:46.92" resultid="16938" heatid="19890" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="216" swimtime="00:00:34.82" resultid="16939" heatid="19949" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="3512" points="141" swimtime="00:03:34.66" resultid="16940" heatid="19994" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5082254" athleteid="17057">
              <RESULTS>
                <RESULT eventid="3547" points="151" swimtime="00:00:50.75" resultid="17058" heatid="19834" lane="2" />
                <RESULT eventid="3590" points="202" swimtime="00:00:40.39" resultid="17060" heatid="19917" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4649975" athleteid="17012">
              <RESULTS>
                <RESULT eventid="3621" points="254" reactiontime="+59" swimtime="00:01:41.76" resultid="17013" heatid="19855" lane="6" entrytime="00:01:42.60" />
                <RESULT eventid="3570" points="260" swimtime="00:02:56.88" resultid="17014" heatid="19873" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="270" reactiontime="+48" swimtime="00:03:36.76" resultid="17015" heatid="19904" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5082249" athleteid="16982">
              <RESULTS>
                <RESULT eventid="3547" points="143" swimtime="00:00:51.66" resultid="16983" heatid="19837" lane="2" entrytime="00:00:47.00" />
                <RESULT eventid="3570" points="135" swimtime="00:03:39.79" resultid="16984" heatid="19875" lane="2" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="161" swimtime="00:00:43.62" resultid="16985" heatid="19920" lane="5" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4489508" athleteid="16402">
              <RESULTS>
                <RESULT eventid="3547" points="230" swimtime="00:00:44.11" resultid="16403" heatid="19838" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="3570" points="233" reactiontime="+81" swimtime="00:03:03.36" resultid="16404" heatid="19873" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="238" swimtime="00:00:38.24" resultid="16405" heatid="19924" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="3505" points="215" swimtime="00:03:28.08" resultid="16406" heatid="19983" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4712853" athleteid="17034">
              <RESULTS>
                <RESULT eventid="3639" points="277" swimtime="00:03:13.45" resultid="17035" heatid="19809" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="307" swimtime="00:00:40.09" resultid="17036" heatid="19839" lane="7" entrytime="00:00:42.50" />
                <RESULT eventid="3570" points="309" reactiontime="+74" swimtime="00:02:47.07" resultid="17037" heatid="19877" lane="3" entrytime="00:02:56.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="326" swimtime="00:00:34.46" resultid="17038" heatid="19926" lane="7" entrytime="00:00:34.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5176269" athleteid="17073">
              <RESULTS>
                <RESULT eventid="3547" points="124" swimtime="00:00:54.14" resultid="17074" heatid="19834" lane="7" />
                <RESULT eventid="3590" points="200" swimtime="00:00:40.52" resultid="17076" heatid="19922" lane="8" entrytime="00:00:40.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4712847" athleteid="17052">
              <RESULTS>
                <RESULT eventid="3639" points="318" swimtime="00:03:04.81" resultid="17053" heatid="19809" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="303" swimtime="00:00:40.28" resultid="17054" heatid="19841" lane="2" entrytime="00:00:37.50" />
                <RESULT eventid="3570" points="313" swimtime="00:02:46.38" resultid="17055" heatid="19879" lane="5" entrytime="00:02:50.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="429" swimtime="00:00:31.44" resultid="17056" heatid="19931" lane="1" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" athleteid="16994">
              <RESULTS>
                <RESULT eventid="3547" points="165" swimtime="00:00:49.27" resultid="16995" heatid="19837" lane="7" entrytime="00:00:47.00" />
                <RESULT comment=" - Start vor dem Startsignal (Zeit: 13:00)" eventid="3570" status="DSQ" swimtime="00:03:40.19" resultid="16996" heatid="19875" lane="3" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="176" swimtime="00:00:42.29" resultid="16997" heatid="19920" lane="4" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" athleteid="16978">
              <RESULTS>
                <RESULT eventid="3547" points="219" swimtime="00:00:44.87" resultid="16979" heatid="19838" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="3570" points="168" swimtime="00:03:24.36" resultid="16980" heatid="19876" lane="1" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="216" swimtime="00:00:39.52" resultid="16981" heatid="19922" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5082247" athleteid="17065">
              <RESULTS>
                <RESULT eventid="3547" points="114" swimtime="00:00:55.78" resultid="17066" heatid="19833" lane="3" />
                <RESULT eventid="3590" points="128" swimtime="00:00:47.07" resultid="17068" heatid="19917" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4902465" athleteid="16941">
              <RESULTS>
                <RESULT eventid="3639" points="262" reactiontime="+73" swimtime="00:03:17.02" resultid="16942" heatid="19812" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="303" swimtime="00:00:40.25" resultid="16943" heatid="19841" lane="6" entrytime="00:00:37.40" />
                <RESULT eventid="3590" points="332" swimtime="00:00:34.26" resultid="16944" heatid="19927" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="3505" points="308" swimtime="00:03:04.77" resultid="16945" heatid="19987" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5093620" athleteid="16990">
              <RESULTS>
                <RESULT eventid="3547" points="127" swimtime="00:00:53.79" resultid="16991" heatid="19837" lane="6" entrytime="00:00:47.00" />
                <RESULT eventid="3570" points="140" swimtime="00:03:37.33" resultid="16992" heatid="19875" lane="6" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="134" swimtime="00:00:46.34" resultid="16993" heatid="19921" lane="8" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5082248" athleteid="17081">
              <RESULTS>
                <RESULT eventid="3547" points="126" swimtime="00:00:53.92" resultid="17082" heatid="19833" lane="6" />
                <RESULT eventid="3590" points="167" swimtime="00:00:43.04" resultid="17084" heatid="19918" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4797141" athleteid="17047">
              <RESULTS>
                <RESULT eventid="3621" points="279" swimtime="00:01:38.56" resultid="17048" heatid="19855" lane="3" entrytime="00:01:42.50" />
                <RESULT eventid="3570" points="276" reactiontime="+65" swimtime="00:02:53.38" resultid="17049" heatid="19874" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="271" reactiontime="+61" swimtime="00:03:36.41" resultid="17050" heatid="19904" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="307" swimtime="00:00:35.15" resultid="17051" heatid="19924" lane="1" entrytime="00:00:36.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4712849" athleteid="17019">
              <RESULTS>
                <RESULT eventid="9711" points="305" reactiontime="+91" swimtime="00:02:49.19" resultid="17020" heatid="19823" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="329" swimtime="00:00:34.79" resultid="17021" heatid="19849" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="3628" points="348" reactiontime="+84" swimtime="00:01:23.26" resultid="17022" heatid="19869" lane="1" entrytime="00:01:24.00" />
                <RESULT eventid="3594" points="381" swimtime="00:00:28.84" resultid="17023" heatid="19953" lane="2" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4104941" athleteid="17002">
              <RESULTS>
                <RESULT eventid="3621" points="270" swimtime="00:01:39.69" resultid="17003" heatid="19856" lane="5" entrytime="00:01:38.50" />
                <RESULT eventid="3570" points="288" reactiontime="+72" swimtime="00:02:51.08" resultid="17004" heatid="19877" lane="6" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="331" swimtime="00:00:34.30" resultid="17005" heatid="19926" lane="4" entrytime="00:00:34.30" />
                <RESULT eventid="3555" points="170" reactiontime="+61" swimtime="00:01:41.04" resultid="17006" heatid="19968" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5164031" athleteid="17077">
              <RESULTS>
                <RESULT eventid="3547" points="116" swimtime="00:00:55.35" resultid="17078" heatid="19833" lane="4" />
                <RESULT eventid="3590" points="110" swimtime="00:00:49.38" resultid="17080" heatid="19917" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4902468" athleteid="16926">
              <RESULTS>
                <RESULT eventid="3551" points="214" swimtime="00:00:40.13" resultid="16927" heatid="19847" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="3649" points="235" swimtime="00:02:45.14" resultid="16928" heatid="19892" lane="5" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="288" swimtime="00:00:31.63" resultid="16929" heatid="19951" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="3562" points="134" reactiontime="+80" swimtime="00:01:37.33" resultid="16930" heatid="19976" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5093618" athleteid="17069">
              <RESULTS>
                <RESULT eventid="3547" points="107" swimtime="00:00:56.86" resultid="17070" heatid="19834" lane="6" />
                <RESULT eventid="3590" points="149" swimtime="00:00:44.74" resultid="17072" heatid="19917" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5164029" athleteid="17061">
              <RESULTS>
                <RESULT eventid="3547" points="161" swimtime="00:00:49.69" resultid="17062" heatid="19833" lane="5" />
                <RESULT eventid="3590" points="194" swimtime="00:00:40.99" resultid="17064" heatid="19921" lane="5" entrytime="00:00:40.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4489509" athleteid="16397">
              <RESULTS>
                <RESULT eventid="3639" points="316" reactiontime="+81" swimtime="00:03:05.16" resultid="16398" heatid="19809" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="275" swimtime="00:00:41.61" resultid="16399" heatid="19839" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="3570" points="341" swimtime="00:02:41.61" resultid="16400" heatid="19878" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="341" swimtime="00:00:33.94" resultid="16401" heatid="19926" lane="3" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4858656" athleteid="17007">
              <RESULTS>
                <RESULT eventid="3547" points="354" swimtime="00:00:38.24" resultid="17008" heatid="19840" lane="1" entrytime="00:00:38.90" />
                <RESULT eventid="3570" points="272" swimtime="00:02:54.33" resultid="17009" heatid="19874" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="274" swimtime="00:00:36.50" resultid="17010" heatid="19925" lane="1" entrytime="00:00:35.50" />
                <RESULT eventid="3505" points="342" swimtime="00:02:58.32" resultid="17011" heatid="19987" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5089299" athleteid="16986">
              <RESULTS>
                <RESULT eventid="3547" points="109" swimtime="00:00:56.60" resultid="16987" heatid="19837" lane="1" entrytime="00:00:47.00" />
                <RESULT eventid="3570" points="119" swimtime="00:03:49.52" resultid="16988" heatid="19875" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="110" swimtime="00:00:49.42" resultid="16989" heatid="19920" lane="2" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5082256" athleteid="16966">
              <RESULTS>
                <RESULT eventid="3621" points="193" swimtime="00:01:51.39" resultid="16967" heatid="19854" lane="5" entrytime="00:01:45.50" />
                <RESULT eventid="3538" points="191" swimtime="00:04:03.20" resultid="16968" heatid="19905" lane="3" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="217" swimtime="00:00:39.44" resultid="16969" heatid="19923" lane="8" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5176268" athleteid="17236">
              <RESULTS>
                <RESULT eventid="3547" points="86" swimtime="00:01:01.29" resultid="17237" heatid="19834" lane="8" />
                <RESULT eventid="3590" points="134" swimtime="00:00:46.29" resultid="17238" heatid="19918" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4649978" athleteid="16931">
              <RESULTS>
                <RESULT eventid="3551" points="126" swimtime="00:00:47.91" resultid="16932" heatid="19847" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="3649" points="164" swimtime="00:03:06.02" resultid="16933" heatid="19890" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="180" swimtime="00:00:37.03" resultid="16934" heatid="19949" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="3562" points="74" swimtime="00:01:58.35" resultid="16935" heatid="19976" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="ITA" swrid="4994490" athleteid="16921">
              <RESULTS>
                <RESULT eventid="3551" points="211" swimtime="00:00:40.33" resultid="16922" heatid="19848" lane="1" entrytime="00:00:41.50" />
                <RESULT eventid="3649" points="214" reactiontime="+76" swimtime="00:02:50.41" resultid="16923" heatid="19892" lane="2" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="233" swimtime="00:00:33.94" resultid="16924" heatid="19950" lane="6" entrytime="00:00:33.40" />
                <RESULT eventid="3512" points="183" swimtime="00:03:16.94" resultid="16925" heatid="19995" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="5089301" athleteid="16970">
              <RESULTS>
                <RESULT eventid="3547" points="140" swimtime="00:00:52.06" resultid="16971" heatid="19838" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="3570" points="203" swimtime="00:03:12.01" resultid="16972" heatid="19876" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="204" swimtime="00:00:40.29" resultid="16973" heatid="19923" lane="7" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="ITA" swrid="4649968" athleteid="17043">
              <RESULTS>
                <RESULT eventid="3621" points="287" reactiontime="+56" swimtime="00:01:37.67" resultid="17044" heatid="19858" lane="4" entrytime="00:01:32.00" />
                <RESULT eventid="3570" points="241" reactiontime="+52" swimtime="00:03:01.34" resultid="17045" heatid="19876" lane="4" entrytime="00:02:59.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="270" reactiontime="+70" swimtime="00:03:36.60" resultid="17046" heatid="19905" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BIEL" nation="SUI" region="RZW" clubid="13007" swrid="65714" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4688265" athleteid="17473">
              <RESULTS>
                <RESULT eventid="3551" points="515" swimtime="00:00:29.99" resultid="17474" heatid="19852" lane="8" entrytime="00:00:29.78" />
                <RESULT eventid="3628" points="461" reactiontime="+74" swimtime="00:01:15.81" resultid="17475" heatid="19872" lane="7" entrytime="00:01:11.07" />
                <RESULT eventid="3594" points="492" swimtime="00:00:26.48" resultid="17476" heatid="19956" lane="1" entrytime="00:00:27.26" />
                <RESULT eventid="3512" points="432" swimtime="00:02:27.94" resultid="17477" heatid="20000" lane="5" entrytime="00:02:21.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="493" swimtime="00:01:05.71" resultid="17478" heatid="20022" lane="7" entrytime="00:01:02.90" />
                <RESULT eventid="3530" points="560" reactiontime="+73" swimtime="00:00:56.89" resultid="17479" heatid="20110" lane="4" entrytime="00:00:57.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4396758" athleteid="17467">
              <RESULTS>
                <RESULT eventid="3649" points="596" reactiontime="+73" swimtime="00:02:01.16" resultid="17468" heatid="19899" lane="6" entrytime="00:01:58.89">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="480" reactiontime="+61" swimtime="00:02:42.58" resultid="17469" heatid="19916" lane="1" entrytime="00:02:36.57">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="521" swimtime="00:00:25.98" resultid="17470" heatid="19958" lane="2" entrytime="00:00:25.88" />
                <RESULT eventid="3519" points="496" swimtime="00:00:33.67" resultid="17471" heatid="20084" lane="8" entrytime="00:00:34.42" />
                <RESULT eventid="3530" points="600" swimtime="00:00:55.61" resultid="17472" heatid="20111" lane="5" entrytime="00:00:55.62" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="5134253" athleteid="17487">
              <RESULTS>
                <RESULT eventid="3594" points="109" swimtime="00:00:43.73" resultid="17488" heatid="19946" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="3519" points="110" swimtime="00:00:55.51" resultid="17489" heatid="20077" lane="5" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="SUI" swrid="4688266" athleteid="17480">
              <RESULTS>
                <RESULT eventid="3551" points="293" swimtime="00:00:36.17" resultid="17481" heatid="19849" lane="7" entrytime="00:00:35.82" />
                <RESULT eventid="3594" points="281" swimtime="00:00:31.92" resultid="17482" heatid="19951" lane="8" entrytime="00:00:32.33" />
                <RESULT eventid="3512" points="295" swimtime="00:02:48.04" resultid="17483" heatid="19998" lane="8" entrytime="00:02:50.02">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="272" swimtime="00:01:20.07" resultid="17484" heatid="20017" lane="3" entrytime="00:01:18.72" />
                <RESULT eventid="3519" points="375" swimtime="00:00:36.96" resultid="17485" heatid="20083" lane="1" entrytime="00:00:37.18" />
                <RESULT eventid="3530" points="295" reactiontime="+62" swimtime="00:01:10.44" resultid="17486" heatid="20105" lane="3" entrytime="00:01:10.02" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="HALL" nation="AUT" region="TLSV" clubid="13734" swrid="68005" name="Breedy Badger">
          <CONTACT city="Innsbruck" email="staatl.t.patrick.holst@gmail.com" name="Breedy Badger" street="Templstrasse" zip="6020" />
          <ATHLETES>
            <ATHLETE birthdate="2003-12-25" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="40037" swrid="4796700" athleteid="17878">
              <RESULTS>
                <RESULT eventid="9711" points="183" reactiontime="+66" swimtime="00:03:20.73" resultid="17879" heatid="19823" lane="3" entrytime="00:03:32.69">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="106" reactiontime="+70" swimtime="00:01:45.23" resultid="17880" heatid="19976" lane="6" />
                <RESULT eventid="3578" points="182" swimtime="00:06:28.21" resultid="17881" heatid="20051" lane="3" entrytime="00:06:24.79">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.14" />
                    <SPLIT distance="200" swimtime="00:03:13.59" />
                    <SPLIT distance="300" swimtime="00:04:53.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="184" swimtime="00:00:46.84" resultid="17882" heatid="20078" lane="2" entrytime="00:00:51.16" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-02-10" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="39895" swrid="4796698" athleteid="17883">
              <RESULTS>
                <RESULT eventid="3621" points="230" swimtime="00:01:45.11" resultid="17884" heatid="19853" lane="2" />
                <RESULT eventid="3555" points="104" reactiontime="+54" swimtime="00:01:58.86" resultid="17885" heatid="19968" lane="7" />
                <RESULT eventid="3598" points="230" swimtime="00:01:34.85" resultid="17886" heatid="20002" lane="3" />
                <RESULT eventid="3523" points="214" swimtime="00:01:26.96" resultid="17887" heatid="20085" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-09-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="43302" swrid="4953379" athleteid="17907">
              <RESULTS>
                <RESULT eventid="3649" points="177" swimtime="00:03:01.62" resultid="17908" heatid="19889" lane="3" entrytime="00:03:15.21">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="188" reactiontime="+91" swimtime="00:03:42.16" resultid="17909" heatid="19911" lane="6" entrytime="00:03:41.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="163" swimtime="00:01:34.97" resultid="17910" heatid="20013" lane="5" entrytime="00:01:37.27" />
                <RESULT eventid="3530" points="196" swimtime="00:01:20.68" resultid="17911" heatid="20101" lane="8" entrytime="00:01:28.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-05-29" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40022" swrid="4796692" athleteid="17992">
              <RESULTS>
                <RESULT eventid="3639" points="263" swimtime="00:03:16.67" resultid="17993" heatid="19811" lane="3" entrytime="00:03:15.18">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="276" swimtime="00:03:11.51" resultid="17994" heatid="19984" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="255" swimtime="00:01:31.63" resultid="17995" heatid="20005" lane="4" entrytime="00:01:27.25" />
                <RESULT eventid="3617" points="230" swimtime="00:00:40.89" resultid="17996" heatid="20025" lane="2" entrytime="00:00:44.09" />
                <RESULT eventid="3523" points="289" swimtime="00:01:18.72" resultid="17997" heatid="20092" lane="8" entrytime="00:01:11.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-11-23" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="40026" swrid="4742493" athleteid="17958">
              <RESULTS>
                <RESULT eventid="3649" points="289" reactiontime="+83" swimtime="00:02:34.25" resultid="17959" heatid="19892" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="261" swimtime="00:00:32.69" resultid="17960" heatid="19950" lane="7" entrytime="00:00:34.26" />
                <RESULT eventid="3512" points="239" swimtime="00:03:00.31" resultid="17961" heatid="19997" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="292" swimtime="00:05:31.68" resultid="17962" heatid="20053" lane="3" entrytime="00:05:53.60">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="200" swimtime="00:02:39.14" />
                    <SPLIT distance="300" swimtime="00:04:06.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="270" reactiontime="+81" swimtime="00:01:12.51" resultid="17963" heatid="20104" lane="6" entrytime="00:01:13.52" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-10-14" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42238" swrid="4992314" athleteid="17924">
              <RESULTS>
                <RESULT eventid="3598" points="238" swimtime="00:01:33.73" resultid="17925" heatid="20003" lane="6" entrytime="00:01:36.49" />
                <RESULT eventid="3514" points="225" swimtime="00:00:48.99" resultid="17926" heatid="20069" lane="3" entrytime="00:00:54.63" />
                <RESULT eventid="3523" points="223" swimtime="00:01:25.74" resultid="17927" heatid="20086" lane="2" entrytime="00:01:28.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-18" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="35095" swrid="4287000" athleteid="17912">
              <RESULTS>
                <RESULT eventid="3639" points="571" reactiontime="+56" swimtime="00:02:32.02" resultid="17913" heatid="19820" lane="4" entrytime="00:02:36.85">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="579" reactiontime="+56" swimtime="00:01:17.32" resultid="17914" heatid="19863" lane="3" entrytime="00:01:15.97" />
                <RESULT eventid="3590" points="625" swimtime="00:00:27.74" resultid="17915" heatid="19937" lane="5" entrytime="00:00:27.49" />
                <RESULT eventid="3617" points="623" swimtime="00:00:29.34" resultid="17916" heatid="20031" lane="5" entrytime="00:00:29.58" />
                <RESULT eventid="3658" points="536" reactiontime="+73" swimtime="00:04:54.31" resultid="17917" heatid="20049" lane="2" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="200" swimtime="00:02:24.00" />
                    <SPLIT distance="300" swimtime="00:03:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="651" swimtime="00:00:34.37" resultid="17918" heatid="20075" lane="4" entrytime="00:00:33.29" />
                <RESULT eventid="15921" points="587" swimtime="00:00:28.33" resultid="20159" heatid="20120" lane="5" late="yes" />
                <RESULT eventid="15972" points="572" swimtime="00:00:28.58" resultid="20160" heatid="20122" lane="5" late="yes" />
                <RESULT eventid="15975" points="565" swimtime="00:00:28.70" resultid="20161" heatid="20124" lane="5" late="yes" />
                <RESULT eventid="15978" points="581" swimtime="00:00:28.43" resultid="20162" heatid="20126" lane="5" late="yes" />
                <RESULT eventid="15981" points="595" swimtime="00:00:28.20" resultid="20163" heatid="20128" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="5172686" athleteid="18458">
              <RESULTS>
                <RESULT eventid="3590" points="166" swimtime="00:00:43.16" resultid="18459" heatid="19918" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-12-04" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41066" swrid="4982373" athleteid="17933">
              <RESULTS>
                <RESULT eventid="3639" points="395" reactiontime="+65" swimtime="00:02:51.82" resultid="17934" heatid="19817" lane="2" entrytime="00:02:50.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="352" reactiontime="+81" swimtime="00:01:31.23" resultid="17935" heatid="19858" lane="6" entrytime="00:01:32.87" />
                <RESULT eventid="3570" points="380" reactiontime="+67" swimtime="00:02:35.92" resultid="17936" heatid="19882" lane="1" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="388" swimtime="00:00:32.51" resultid="17937" heatid="19929" lane="6" entrytime="00:00:32.13" />
                <RESULT eventid="3598" points="319" swimtime="00:01:25.06" resultid="17938" heatid="20005" lane="6" entrytime="00:01:27.70" />
                <RESULT eventid="3658" points="371" swimtime="00:05:32.57" resultid="17939" heatid="20047" lane="3" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="200" swimtime="00:02:42.42" />
                    <SPLIT distance="300" swimtime="00:04:08.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-05-10" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40030" swrid="4796693" athleteid="17919">
              <RESULTS>
                <RESULT eventid="3639" points="226" reactiontime="+72" swimtime="00:03:26.81" resultid="17920" heatid="19809" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="289" swimtime="00:00:35.89" resultid="17921" heatid="19922" lane="5" entrytime="00:00:39.25" />
                <RESULT eventid="3658" points="205" reactiontime="+65" swimtime="00:06:44.97" resultid="17922" heatid="20040" lane="3" entrytime="00:08:12.76">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.50" />
                    <SPLIT distance="200" swimtime="00:03:16.61" />
                    <SPLIT distance="300" swimtime="00:05:03.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="249" swimtime="00:00:47.35" resultid="17923" heatid="20070" lane="7" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="5190735" athleteid="17975">
              <RESULTS>
                <RESULT comment=" - Start vor dem Startsignal (Zeit: 12:52)" eventid="3570" status="DSQ" swimtime="00:03:22.89" resultid="17976" heatid="19873" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="185" swimtime="00:04:05.75" resultid="17977" heatid="19905" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3617" points="157" swimtime="00:00:46.40" resultid="17978" heatid="20023" lane="6" />
                <RESULT eventid="3523" points="162" reactiontime="+84" swimtime="00:01:35.51" resultid="17979" heatid="20085" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-13" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="31928" swrid="4078016" athleteid="17888">
              <RESULTS>
                <RESULT eventid="3639" points="593" reactiontime="+62" swimtime="00:02:30.11" resultid="17889" heatid="19822" lane="7" entrytime="00:02:30.19">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="609" reactiontime="+56" swimtime="00:02:13.27" resultid="17890" heatid="19888" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="543" swimtime="00:00:29.07" resultid="17891" heatid="19937" lane="1" entrytime="00:00:29.09" />
                <RESULT eventid="3555" points="563" reactiontime="+61" swimtime="00:01:07.89" resultid="17892" heatid="19975" lane="8" entrytime="00:01:08.50" />
                <RESULT eventid="3658" points="609" reactiontime="+70" swimtime="00:04:42.06" resultid="17893" heatid="20049" lane="7" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="200" swimtime="00:02:18.80" />
                    <SPLIT distance="300" swimtime="00:03:30.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-03-07" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="42771" swrid="5071977" athleteid="17872">
              <RESULTS>
                <RESULT eventid="3551" points="222" swimtime="00:00:39.65" resultid="17873" heatid="19846" lane="3" entrytime="00:00:46.48" />
                <RESULT eventid="3649" points="192" reactiontime="+52" swimtime="00:02:56.65" resultid="17874" heatid="19890" lane="8" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="236" swimtime="00:03:00.94" resultid="17875" heatid="19995" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="224" swimtime="00:01:25.45" resultid="17876" heatid="20016" lane="7" entrytime="00:01:25.00" />
                <RESULT eventid="3530" points="207" reactiontime="+54" swimtime="00:01:19.30" resultid="17877" heatid="20102" lane="8" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-11-23" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="37027" swrid="4478903" athleteid="17855">
              <RESULTS>
                <RESULT eventid="9711" points="449" reactiontime="+71" swimtime="00:02:28.77" resultid="17856" heatid="19830" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="444" swimtime="00:02:13.61" resultid="17857" heatid="19897" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="473" reactiontime="+71" swimtime="00:01:03.92" resultid="17858" heatid="19980" lane="5" entrytime="00:01:04.00" />
                <RESULT eventid="3613" points="500" swimtime="00:00:28.25" resultid="17859" heatid="20038" lane="3" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-06-03" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="40035" swrid="4796701" athleteid="17900">
              <RESULTS>
                <RESULT eventid="9711" points="279" swimtime="00:02:54.33" resultid="17901" heatid="19825" lane="5" entrytime="00:03:03.99">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="298" reactiontime="+88" swimtime="00:01:27.61" resultid="17902" heatid="19866" lane="4" entrytime="00:01:32.13" />
                <RESULT eventid="3545" points="273" reactiontime="+79" swimtime="00:03:16.20" resultid="17903" heatid="19912" lane="2" entrytime="00:03:26.29">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="226" swimtime="00:01:25.17" resultid="17904" heatid="20015" lane="6" entrytime="00:01:27.20" />
                <RESULT eventid="3578" points="248" reactiontime="+78" swimtime="00:05:50.23" resultid="17905" heatid="20054" lane="1" entrytime="00:05:39.95">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.42" />
                    <SPLIT distance="200" swimtime="00:02:49.32" />
                    <SPLIT distance="300" swimtime="00:04:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="324" reactiontime="+82" swimtime="00:01:08.27" resultid="17906" heatid="20105" lane="7" entrytime="00:01:11.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-12-28" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="43300" swrid="4953380" athleteid="17980">
              <RESULTS>
                <RESULT eventid="3551" points="202" swimtime="00:00:40.92" resultid="17981" heatid="19847" lane="3" entrytime="00:00:42.10" />
                <RESULT eventid="3649" points="244" reactiontime="+83" swimtime="00:02:43.06" resultid="17982" heatid="19892" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="211" swimtime="00:03:07.72" resultid="17983" heatid="19997" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="198" swimtime="00:01:28.98" resultid="17984" heatid="20016" lane="2" entrytime="00:01:25.00" />
                <RESULT eventid="3578" points="251" reactiontime="+83" swimtime="00:05:48.44" resultid="17985" heatid="20051" lane="4" entrytime="00:06:18.18">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.42" />
                    <SPLIT distance="200" swimtime="00:02:52.08" />
                    <SPLIT distance="300" swimtime="00:04:22.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-09-05" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="5172683" athleteid="17967">
              <RESULTS>
                <RESULT eventid="3551" points="51" swimtime="00:01:04.77" resultid="17968" heatid="19845" lane="5" />
                <RESULT eventid="3594" points="57" swimtime="00:00:54.23" resultid="17969" heatid="19945" lane="4" />
                <RESULT comment=" - Start vor dem Startsignal (Zeit: 13:56)" eventid="3519" status="DSQ" swimtime="00:01:05.02" resultid="17970" heatid="20076" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-02-04" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="37566" swrid="4487226" athleteid="17865">
              <RESULTS>
                <RESULT eventid="9711" points="414" reactiontime="+69" swimtime="00:02:32.90" resultid="17866" heatid="19831" lane="1" entrytime="00:02:26.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="406" swimtime="00:00:32.45" resultid="17867" heatid="19851" lane="2" entrytime="00:00:30.96" />
                <RESULT eventid="3594" points="413" swimtime="00:00:28.07" resultid="17868" heatid="19952" lane="7" entrytime="00:00:30.36" />
                <RESULT eventid="3512" points="449" swimtime="00:02:26.06" resultid="17869" heatid="20000" lane="2" entrytime="00:02:23.63">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="445" swimtime="00:01:08.02" resultid="17870" heatid="20021" lane="8" entrytime="00:01:07.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-06-05" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42237" swrid="4992315" athleteid="17928">
              <RESULTS>
                <RESULT eventid="3547" points="270" swimtime="00:00:41.86" resultid="17929" heatid="19838" lane="2" entrytime="00:00:44.41" />
                <RESULT eventid="3590" points="342" swimtime="00:00:33.93" resultid="17930" heatid="19924" lane="7" entrytime="00:00:36.37" />
                <RESULT eventid="3617" points="265" swimtime="00:00:39.02" resultid="17931" heatid="20026" lane="8" entrytime="00:00:41.58" />
                <RESULT eventid="3514" points="246" swimtime="00:00:47.50" resultid="17932" heatid="20070" lane="2" entrytime="00:00:51.06" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-08-10" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="40021" swrid="4796690" athleteid="17998">
              <RESULTS>
                <RESULT eventid="9711" points="279" reactiontime="+60" swimtime="00:02:54.31" resultid="17999" heatid="19827" lane="7" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="269" reactiontime="+73" swimtime="00:01:30.74" resultid="18000" heatid="19867" lane="7" entrytime="00:01:31.03" />
                <RESULT eventid="3605" points="274" swimtime="00:01:19.91" resultid="18002" heatid="20017" lane="7" entrytime="00:01:20.81" />
                <RESULT eventid="3530" points="312" reactiontime="+65" swimtime="00:01:09.15" resultid="18003" heatid="20105" lane="8" entrytime="00:01:11.74" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-11-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="38064" swrid="4932701" athleteid="17947">
              <RESULTS>
                <RESULT eventid="9711" points="170" reactiontime="+78" swimtime="00:03:25.40" resultid="17948" heatid="19823" lane="6" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="136" reactiontime="+67" swimtime="00:03:17.99" resultid="17949" heatid="19889" lane="6" entrytime="00:03:19.62">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="166" swimtime="00:03:51.20" resultid="17950" heatid="19911" lane="2" entrytime="00:03:49.13">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="144" swimtime="00:03:33.36" resultid="17951" heatid="19994" lane="5" entrytime="00:03:25.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-10-24" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="40393" swrid="4796702" athleteid="17952">
              <RESULTS>
                <RESULT eventid="9711" points="241" reactiontime="+68" swimtime="00:03:03.14" resultid="17953" heatid="19826" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="305" swimtime="00:01:27.00" resultid="17954" heatid="19867" lane="3" entrytime="00:01:30.00" />
                <RESULT eventid="3545" points="307" swimtime="00:03:08.64" resultid="17955" heatid="19913" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="206" swimtime="00:03:09.35" resultid="17956" heatid="19996" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="328" swimtime="00:00:38.67" resultid="17957" heatid="20080" lane="6" entrytime="00:00:42.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-11-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="4932694" athleteid="17860">
              <RESULTS>
                <RESULT eventid="3621" points="141" swimtime="00:02:03.78" resultid="17861" heatid="19853" lane="6" />
                <RESULT eventid="3505" points="154" swimtime="00:03:52.82" resultid="17862" heatid="19983" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" status="DNS" swimtime="00:00:00.00" resultid="17863" heatid="20002" lane="5" />
                <RESULT eventid="3523" points="136" swimtime="00:01:41.21" resultid="17864" heatid="20085" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-10-18" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="37266" swrid="4639766" athleteid="17964">
              <RESULTS>
                <RESULT eventid="3578" points="549" reactiontime="+47" swimtime="00:04:28.73" resultid="17965" heatid="20058" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.19" />
                    <SPLIT distance="200" swimtime="00:02:07.23" />
                    <SPLIT distance="300" swimtime="00:03:18.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="527" reactiontime="+74" swimtime="00:05:01.83" resultid="17966" heatid="20119" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="200" swimtime="00:02:27.48" />
                    <SPLIT distance="300" swimtime="00:03:53.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-02-11" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="37563" swrid="4656765" athleteid="17940">
              <RESULTS>
                <RESULT eventid="3570" points="510" swimtime="00:02:21.39" resultid="17941" heatid="19887" lane="5" entrytime="00:02:14.86">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="526" swimtime="00:00:29.38" resultid="17942" heatid="19937" lane="7" entrytime="00:00:28.87" />
                <RESULT eventid="3617" points="545" swimtime="00:00:30.68" resultid="17943" heatid="20030" lane="3" entrytime="00:00:31.58" />
                <RESULT eventid="3523" points="556" reactiontime="+60" swimtime="00:01:03.29" resultid="17944" heatid="20098" lane="3" entrytime="00:01:03.31" />
                <RESULT eventid="3639" points="463" swimtime="00:02:43.04" resultid="17945" heatid="19820" lane="5" entrytime="00:02:36.97">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3636" points="504" reactiontime="+65" swimtime="00:05:38.49" resultid="17946" heatid="20115" lane="5" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="200" swimtime="00:02:40.06" />
                    <SPLIT distance="300" swimtime="00:04:20.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-04-14" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42236" swrid="4992316" athleteid="17986">
              <RESULTS>
                <RESULT eventid="3639" points="289" swimtime="00:03:10.76" resultid="17987" heatid="19809" lane="4" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="259" swimtime="00:03:39.78" resultid="17988" heatid="19906" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="210" swimtime="00:01:34.17" resultid="17989" heatid="19969" lane="4" entrytime="00:01:30.00" />
                <RESULT eventid="3617" points="307" swimtime="00:00:37.16" resultid="17990" heatid="20026" lane="6" entrytime="00:00:40.48" />
                <RESULT eventid="3586" points="211" swimtime="00:03:24.42" resultid="17991" heatid="20063" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-04-21" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40036" swrid="4796688" athleteid="17894">
              <RESULTS>
                <RESULT eventid="3639" points="310" swimtime="00:03:06.22" resultid="17895" heatid="19811" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="367" reactiontime="+88" swimtime="00:01:30.00" resultid="17896" heatid="19859" lane="2" entrytime="00:01:30.00" />
                <RESULT eventid="3538" points="367" swimtime="00:03:15.64" resultid="17897" heatid="19907" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3658" points="270" reactiontime="+68" swimtime="00:06:09.65" resultid="17898" heatid="20041" lane="2" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.41" />
                    <SPLIT distance="200" swimtime="00:03:03.64" />
                    <SPLIT distance="300" swimtime="00:04:40.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="381" swimtime="00:00:41.09" resultid="17899" heatid="20071" lane="3" entrytime="00:00:45.04" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-10-18" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="5172684" athleteid="17971">
              <RESULTS>
                <RESULT eventid="3551" points="19" swimtime="00:01:29.87" resultid="17972" heatid="19845" lane="3" />
                <RESULT eventid="3594" points="10" swimtime="00:01:34.97" resultid="17973" heatid="19945" lane="5" />
                <RESULT eventid="3519" points="57" swimtime="00:01:08.93" resultid="17974" heatid="20076" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SUGS" nation="AUT" region="SLSV" clubid="13021" swrid="65818" name="Breedy Badger">
          <CONTACT email="hanni.gerstbauer@gmx.at" name="Breedy Badger" />
          <ATHLETES>
            <ATHLETE birthdate="2004-09-08" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="5101399" athleteid="16879">
              <RESULTS>
                <RESULT eventid="9711" points="229" swimtime="00:03:06.22" resultid="17281" heatid="19824" lane="3" entrytime="00:03:17.75">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="246" swimtime="00:02:42.72" resultid="17282" heatid="19890" lane="3" entrytime="00:02:51.67">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="202" swimtime="00:03:10.55" resultid="17283" heatid="19995" lane="3" entrytime="00:03:10.98">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="176" swimtime="00:01:32.68" resultid="17284" heatid="20014" lane="2" entrytime="00:01:32.45" />
                <RESULT eventid="3578" points="279" reactiontime="+72" swimtime="00:05:36.52" resultid="17285" heatid="20052" lane="2" entrytime="00:06:02.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.25" />
                    <SPLIT distance="200" swimtime="00:02:47.45" />
                    <SPLIT distance="300" swimtime="00:04:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="236" swimtime="00:01:15.84" resultid="17286" heatid="20101" lane="5" entrytime="00:01:20.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-05-21" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="4841398" athleteid="16900">
              <RESULTS>
                <RESULT eventid="9711" points="233" swimtime="00:03:05.03" resultid="17299" heatid="19825" lane="2" entrytime="00:03:12.43">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="249" swimtime="00:02:42.13" resultid="17300" heatid="19891" lane="2" entrytime="00:02:48.67">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="237" swimtime="00:03:00.78" resultid="17301" heatid="19996" lane="5" entrytime="00:03:00.12">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="214" swimtime="00:01:26.75" resultid="17302" heatid="20015" lane="5" entrytime="00:01:26.45" />
                <RESULT comment=" - Start vor dem Startsignal (Zeit: 11:56)" eventid="3578" status="DSQ" swimtime="00:05:36.04" resultid="17303" heatid="20053" lane="8" entrytime="00:05:59.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.80" />
                    <SPLIT distance="200" swimtime="00:02:41.30" />
                    <SPLIT distance="300" swimtime="00:04:08.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="234" reactiontime="+63" swimtime="00:01:16.02" resultid="17304" heatid="20102" lane="7" entrytime="00:01:19.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-09-13" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="4895337" athleteid="16886">
              <RESULTS>
                <RESULT eventid="9711" points="243" swimtime="00:03:02.45" resultid="17287" heatid="19825" lane="1" entrytime="00:03:12.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="269" swimtime="00:02:37.84" resultid="17288" heatid="19891" lane="8" entrytime="00:02:49.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="234" swimtime="00:03:01.51" resultid="17289" heatid="19996" lane="6" entrytime="00:03:01.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="210" swimtime="00:01:27.38" resultid="17290" heatid="20015" lane="8" entrytime="00:01:29.54" />
                <RESULT eventid="3578" points="284" swimtime="00:05:34.56" resultid="17291" heatid="20052" lane="6" entrytime="00:06:02.08">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                    <SPLIT distance="200" swimtime="00:02:46.03" />
                    <SPLIT distance="300" swimtime="00:04:12.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="271" swimtime="00:01:12.48" resultid="17292" heatid="20102" lane="5" entrytime="00:01:18.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-02-12" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" swrid="4789286" athleteid="16893">
              <RESULTS>
                <RESULT eventid="3628" points="315" swimtime="00:01:26.08" resultid="17293" heatid="19867" lane="4" entrytime="00:01:27.59" />
                <RESULT eventid="3649" points="281" swimtime="00:02:35.57" resultid="17294" heatid="19891" lane="3" entrytime="00:02:48.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="319" reactiontime="+52" swimtime="00:03:06.19" resultid="17295" heatid="19914" lane="8" entrytime="00:03:06.84">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="272" swimtime="00:02:52.53" resultid="17296" heatid="19997" lane="1" entrytime="00:02:59.78">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="292" reactiontime="+47" swimtime="00:05:31.50" resultid="17297" heatid="20053" lane="7" entrytime="00:05:56.78">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                    <SPLIT distance="200" swimtime="00:02:42.68" />
                    <SPLIT distance="300" swimtime="00:04:08.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="293" swimtime="00:00:40.15" resultid="17298" heatid="20081" lane="8" entrytime="00:00:40.72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-03-14" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="4794749" athleteid="16914">
              <RESULTS>
                <RESULT eventid="3639" points="300" reactiontime="+85" swimtime="00:03:08.37" resultid="17311" heatid="19811" lane="8" entrytime="00:03:17.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="292" swimtime="00:02:50.17" resultid="17312" heatid="19877" lane="1" entrytime="00:02:58.97">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="317" swimtime="00:03:03.04" resultid="17313" heatid="19985" lane="4" entrytime="00:03:08.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="302" swimtime="00:01:26.58" resultid="17314" heatid="20005" lane="8" entrytime="00:01:28.78" />
                <RESULT eventid="3658" points="295" swimtime="00:05:59.11" resultid="17315" heatid="20041" lane="4" entrytime="00:06:10.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.47" />
                    <SPLIT distance="200" swimtime="00:02:55.08" />
                    <SPLIT distance="300" swimtime="00:04:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="298" swimtime="00:01:17.91" resultid="17316" heatid="20087" lane="4" entrytime="00:01:19.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-05-13" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" swrid="5001672" athleteid="16907">
              <RESULTS>
                <RESULT eventid="3639" points="307" reactiontime="+66" swimtime="00:03:06.89" resultid="17305" heatid="19812" lane="7" entrytime="00:03:12.45">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="360" swimtime="00:02:38.72" resultid="17306" heatid="19877" lane="5" entrytime="00:02:56.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="339" swimtime="00:02:58.92" resultid="17307" heatid="19986" lane="2" entrytime="00:03:05.78">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="320" swimtime="00:01:24.89" resultid="17308" heatid="20005" lane="1" entrytime="00:01:28.50" />
                <RESULT eventid="3658" points="349" swimtime="00:05:39.62" resultid="17309" heatid="20043" lane="5" entrytime="00:05:52.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="200" swimtime="00:02:45.35" />
                    <SPLIT distance="300" swimtime="00:04:14.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="362" reactiontime="+49" swimtime="00:01:13.03" resultid="17310" heatid="20089" lane="4" entrytime="00:01:15.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AUGSB" nation="GER" region="02" clubid="17317" name="Breedy Badger" shortname="SV Augsburg ">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="264119" swrid="4491214" athleteid="17341">
              <RESULTS>
                <RESULT eventid="3639" points="321" reactiontime="+97" swimtime="00:03:04.05" resultid="17342" heatid="19817" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="407" reactiontime="+84" swimtime="00:02:32.38" resultid="17343" heatid="19885" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="449" swimtime="00:00:30.97" resultid="17344" heatid="19934" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="3505" points="329" swimtime="00:03:00.66" resultid="17345" heatid="19989" lane="6" entrytime="00:02:48.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3617" points="397" swimtime="00:00:34.09" resultid="17346" heatid="20028" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="3523" points="457" swimtime="00:01:07.56" resultid="17347" heatid="20098" lane="5" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="350186" swrid="5063091" athleteid="17366">
              <RESULTS>
                <RESULT eventid="9711" points="250" reactiontime="+65" swimtime="00:03:00.73" resultid="17367" heatid="19827" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="332" reactiontime="+57" swimtime="00:01:24.58" resultid="17368" heatid="19870" lane="3" entrytime="00:01:19.80" />
                <RESULT eventid="3545" points="300" reactiontime="+66" swimtime="00:03:10.04" resultid="17369" heatid="19914" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="341" swimtime="00:00:38.15" resultid="17370" heatid="20083" lane="7" entrytime="00:00:37.10" />
                <RESULT eventid="3530" points="253" reactiontime="+63" swimtime="00:01:14.08" resultid="17371" heatid="20105" lane="6" entrytime="00:01:10.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="310494" swrid="5097997" athleteid="17357">
              <RESULTS>
                <RESULT eventid="9711" points="225" swimtime="00:03:07.16" resultid="17358" heatid="19826" lane="4" entrytime="00:02:58.60">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="176" swimtime="00:00:42.83" resultid="17359" heatid="19848" lane="6" entrytime="00:00:38.60" />
                <RESULT eventid="3649" points="251" reactiontime="+64" swimtime="00:02:41.56" resultid="17360" heatid="19892" lane="7" entrytime="00:02:42.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="238" swimtime="00:00:33.70" resultid="17361" heatid="19950" lane="5" entrytime="00:00:32.80" />
                <RESULT eventid="3512" points="210" swimtime="00:03:08.27" resultid="17362" heatid="19997" lane="6" entrytime="00:02:56.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="192" swimtime="00:01:29.88" resultid="17363" heatid="20016" lane="3" entrytime="00:01:24.30" />
                <RESULT eventid="3613" points="193" swimtime="00:00:38.76" resultid="17364" heatid="20034" lane="6" entrytime="00:00:37.50" />
                <RESULT eventid="3530" points="238" swimtime="00:01:15.61" resultid="17365" heatid="20103" lane="5" entrytime="00:01:15.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="333282" swrid="4973167" athleteid="17348">
              <RESULTS>
                <RESULT eventid="9711" points="355" reactiontime="+55" swimtime="00:02:40.89" resultid="17349" heatid="19828" lane="4" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="370" reactiontime="+55" swimtime="00:02:22.00" resultid="17350" heatid="19894" lane="2" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="433" swimtime="00:00:27.62" resultid="17351" heatid="19959" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="3512" points="332" swimtime="00:02:41.53" resultid="17352" heatid="19998" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="347" swimtime="00:01:13.91" resultid="17353" heatid="20019" lane="6" entrytime="00:01:13.00" />
                <RESULT eventid="3613" points="372" swimtime="00:00:31.18" resultid="17354" heatid="20037" lane="3" entrytime="00:00:30.10" />
                <RESULT eventid="3519" points="329" swimtime="00:00:38.60" resultid="17355" heatid="20083" lane="6" entrytime="00:00:36.20" />
                <RESULT eventid="3530" points="425" reactiontime="+57" swimtime="00:01:02.37" resultid="17356" heatid="20108" lane="4" entrytime="00:01:01.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="186316" swrid="4154164" athleteid="17331">
              <RESULTS>
                <RESULT eventid="9711" points="348" reactiontime="+78" swimtime="00:02:42.07" resultid="17332" heatid="19829" lane="6" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="374" swimtime="00:00:33.36" resultid="17333" heatid="19851" lane="6" entrytime="00:00:30.80" />
                <RESULT eventid="3649" points="365" reactiontime="+78" swimtime="00:02:22.63" resultid="17334" heatid="19895" lane="3" entrytime="00:02:16.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="435" swimtime="00:00:27.59" resultid="17335" heatid="19959" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="3562" points="300" reactiontime="+75" swimtime="00:01:14.36" resultid="17336" heatid="19978" lane="5" entrytime="00:01:11.00" />
                <RESULT eventid="3512" status="DNS" swimtime="00:00:00.00" resultid="17337" heatid="19999" lane="2" entrytime="00:02:34.20" />
                <RESULT eventid="3605" points="366" swimtime="00:01:12.58" resultid="17338" heatid="20020" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="3613" points="385" swimtime="00:00:30.81" resultid="17339" heatid="20038" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="3530" points="433" reactiontime="+74" swimtime="00:01:01.98" resultid="17340" heatid="20110" lane="1" entrytime="00:00:59.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="159017" swrid="4089861" athleteid="17323">
              <RESULTS>
                <RESULT eventid="9711" points="336" swimtime="00:02:43.97" resultid="17324" heatid="19827" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="283" reactiontime="+87" swimtime="00:01:29.20" resultid="17325" heatid="19869" lane="8" entrytime="00:01:24.00" />
                <RESULT eventid="3649" points="350" reactiontime="+87" swimtime="00:02:24.64" resultid="17326" heatid="19894" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="387" swimtime="00:00:28.69" resultid="17327" heatid="19954" lane="4" entrytime="00:00:27.90" />
                <RESULT eventid="3613" points="378" swimtime="00:00:31.01" resultid="17328" heatid="20037" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="3519" points="316" swimtime="00:00:39.14" resultid="17329" heatid="20082" lane="3" entrytime="00:00:37.90" />
                <RESULT eventid="3530" points="413" reactiontime="+81" swimtime="00:01:02.99" resultid="17330" heatid="20109" lane="5" entrytime="00:00:59.70" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OTTOBR" nation="GER" region="02" clubid="16490" name="Breedy Badger" shortname="SV Ottobrunn ">
          <CONTACT city="München-Trudering" email="dirk.opavsky@sv-ottobrunn.de" name="Breedy Badger" phone="+49 171/8153369" street="Hoferichterweg 19a" zip="81827" />
          <ATHLETES>
            <ATHLETE birthdate="2004-06-18" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="345304" swrid="5022160" athleteid="16534">
              <RESULTS>
                <RESULT eventid="3547" points="225" swimtime="00:00:44.47" resultid="18689" heatid="19839" lane="8" entrytime="00:00:42.90" />
                <RESULT eventid="3621" points="239" swimtime="00:01:43.80" resultid="18690" heatid="19856" lane="7" entrytime="00:01:40.72" />
                <RESULT eventid="3538" points="264" swimtime="00:03:38.41" resultid="18691" heatid="19905" lane="6" entrytime="00:03:38.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="255" swimtime="00:03:16.79" resultid="18692" heatid="19985" lane="7" entrytime="00:03:11.26">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="248" swimtime="00:01:32.45" resultid="18693" heatid="20004" lane="3" entrytime="00:01:31.46" />
                <RESULT eventid="3617" points="154" swimtime="00:00:46.76" resultid="18694" heatid="20025" lane="8" entrytime="00:00:45.81" />
                <RESULT eventid="3514" points="268" swimtime="00:00:46.20" resultid="18695" heatid="20071" lane="6" entrytime="00:00:45.41" />
                <RESULT eventid="3523" points="201" swimtime="00:01:28.83" resultid="18696" heatid="20086" lane="7" entrytime="00:01:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-04-15" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="345309" swrid="4973236" athleteid="16520">
              <RESULTS>
                <RESULT eventid="3547" points="275" swimtime="00:00:41.60" resultid="18677" heatid="19839" lane="5" entrytime="00:00:40.87" />
                <RESULT eventid="3621" points="186" swimtime="00:01:52.89" resultid="18678" heatid="19854" lane="8" entrytime="00:01:50.48" />
                <RESULT eventid="3590" points="201" swimtime="00:00:40.48" resultid="18679" heatid="19921" lane="3" entrytime="00:00:40.90" />
                <RESULT eventid="3505" points="253" swimtime="00:03:17.28" resultid="18680" heatid="19984" lane="3" entrytime="00:03:15.43">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="238" swimtime="00:01:33.71" resultid="18681" heatid="20004" lane="2" entrytime="00:01:32.45" />
                <RESULT eventid="3617" points="133" swimtime="00:00:49.07" resultid="18682" heatid="20024" lane="2" entrytime="00:00:49.50" />
                <RESULT eventid="3514" points="195" swimtime="00:00:51.36" resultid="18683" heatid="20070" lane="6" entrytime="00:00:50.82" />
                <RESULT eventid="3523" points="176" swimtime="00:01:32.74" resultid="18684" heatid="20086" lane="1" entrytime="00:01:30.07" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-06-28" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="345302" swrid="4973240" athleteid="16543">
              <RESULTS>
                <RESULT eventid="3639" points="270" swimtime="00:03:14.94" resultid="18697" heatid="19811" lane="2" entrytime="00:03:15.68">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="312" swimtime="00:01:34.95" resultid="18698" heatid="19858" lane="8" entrytime="00:01:34.45" />
                <RESULT eventid="3538" points="310" swimtime="00:03:27.03" resultid="18699" heatid="19906" lane="3" entrytime="00:03:28.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="288" swimtime="00:03:08.97" resultid="18700" heatid="19986" lane="7" entrytime="00:03:06.94">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="289" swimtime="00:01:27.89" resultid="18701" heatid="20005" lane="5" entrytime="00:01:27.51" />
                <RESULT eventid="3617" points="192" swimtime="00:00:43.39" resultid="18702" heatid="20025" lane="6" entrytime="00:00:42.96" />
                <RESULT eventid="3514" points="347" swimtime="00:00:42.38" resultid="18703" heatid="20072" lane="8" entrytime="00:00:44.75" />
                <RESULT eventid="3523" points="223" swimtime="00:01:25.83" resultid="18704" heatid="20086" lane="3" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-10-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="345300" swrid="4973242" athleteid="16561">
              <RESULTS>
                <RESULT eventid="3551" points="238" swimtime="00:00:38.76" resultid="18713" heatid="19848" lane="4" entrytime="00:00:36.45" />
                <RESULT eventid="3649" points="211" reactiontime="+68" swimtime="00:02:51.13" resultid="18714" heatid="19891" lane="1" entrytime="00:02:49.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="173" reactiontime="+63" swimtime="00:03:48.16" resultid="18715" heatid="19912" lane="7" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="233" swimtime="00:03:01.68" resultid="18716" heatid="19997" lane="3" entrytime="00:02:55.92">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="243" swimtime="00:01:23.19" resultid="18717" heatid="20016" lane="4" entrytime="00:01:22.30" />
                <RESULT eventid="3578" points="197" swimtime="00:06:18.17" resultid="18718" heatid="20053" lane="2" entrytime="00:05:54.85">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.10" />
                    <SPLIT distance="200" swimtime="00:03:03.48" />
                    <SPLIT distance="300" swimtime="00:04:41.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-04-07" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="345310" swrid="4973235" athleteid="16511">
              <RESULTS>
                <RESULT eventid="9711" points="219" swimtime="00:03:08.90" resultid="18669" heatid="19824" lane="5" entrytime="00:03:17.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="181" swimtime="00:01:43.37" resultid="18670" heatid="19864" lane="5" entrytime="00:01:45.00" />
                <RESULT eventid="3545" points="178" swimtime="00:03:46.04" resultid="18671" heatid="19911" lane="3" entrytime="00:03:41.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="246" swimtime="00:00:33.36" resultid="18672" heatid="19950" lane="1" entrytime="00:00:34.44" />
                <RESULT eventid="3605" points="209" swimtime="00:01:27.48" resultid="18673" heatid="20015" lane="3" entrytime="00:01:26.55" />
                <RESULT eventid="3578" points="236" swimtime="00:05:55.73" resultid="18674" heatid="20051" lane="5" entrytime="00:06:21.69">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="200" swimtime="00:02:55.79" />
                    <SPLIT distance="300" swimtime="00:04:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="174" swimtime="00:00:47.76" resultid="18675" heatid="20078" lane="3" entrytime="00:00:50.64" />
                <RESULT eventid="3530" points="274" reactiontime="+68" swimtime="00:01:12.18" resultid="18676" heatid="20103" lane="7" entrytime="00:01:17.07" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-06-12" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="380866" athleteid="16502">
              <RESULTS>
                <RESULT comment=" - Anschlag nicht in Rückenlage (Zeit: 11:19)" eventid="9711" status="DSQ" swimtime="00:03:28.07" resultid="18661" heatid="19823" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="199" reactiontime="+57" swimtime="00:01:40.26" resultid="18662" heatid="19865" lane="1" entrytime="00:01:38.64" />
                <RESULT eventid="3545" points="218" reactiontime="+52" swimtime="00:03:31.48" resultid="18663" heatid="19912" lane="1" entrytime="00:03:29.05">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="166" swimtime="00:03:23.48" resultid="18664" heatid="19994" lane="3" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="151" swimtime="00:01:37.33" resultid="18665" heatid="20014" lane="8" entrytime="00:01:35.72" />
                <RESULT eventid="3613" points="86" swimtime="00:00:50.77" resultid="18666" heatid="20033" lane="8" entrytime="00:00:50.00" />
                <RESULT eventid="3519" points="208" swimtime="00:00:44.98" resultid="18667" heatid="20079" lane="3" entrytime="00:00:46.63" />
                <RESULT eventid="3530" points="154" reactiontime="+48" swimtime="00:01:27.41" resultid="18668" heatid="20101" lane="2" entrytime="00:01:24.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="362017" swrid="5066101" athleteid="16552">
              <RESULTS>
                <RESULT eventid="3639" points="230" swimtime="00:03:25.77" resultid="18705" heatid="19810" lane="5" entrytime="00:03:20.81">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="258" swimtime="00:00:42.47" resultid="18706" heatid="19840" lane="7" entrytime="00:00:38.83" />
                <RESULT eventid="3570" points="235" swimtime="00:03:03.04" resultid="18707" heatid="19877" lane="8" entrytime="00:02:59.89">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="297" swimtime="00:00:35.53" resultid="18708" heatid="19926" lane="1" entrytime="00:00:34.89" />
                <RESULT eventid="3505" points="265" swimtime="00:03:14.30" resultid="18709" heatid="19985" lane="2" entrytime="00:03:10.47">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="258" swimtime="00:01:31.28" resultid="18710" heatid="20004" lane="4" entrytime="00:01:29.08" />
                <RESULT eventid="3658" points="218" swimtime="00:06:36.78" resultid="18711" heatid="20040" lane="5" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                    <SPLIT distance="200" swimtime="00:03:12.81" />
                    <SPLIT distance="300" swimtime="00:04:57.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="277" swimtime="00:01:19.85" resultid="18712" heatid="20088" lane="2" entrytime="00:01:17.86" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-09-04" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="345299" swrid="4973239" athleteid="16568">
              <RESULTS>
                <RESULT eventid="3547" status="DNS" swimtime="00:00:00.00" resultid="18719" heatid="19841" lane="8" entrytime="00:00:37.75" />
                <RESULT eventid="3621" status="DNS" swimtime="00:00:00.00" resultid="18720" heatid="19855" lane="4" entrytime="00:01:41.35" />
                <RESULT eventid="3555" status="DNS" swimtime="00:00:00.00" resultid="18721" heatid="19969" lane="8" entrytime="00:01:35.07" />
                <RESULT eventid="3505" status="DNS" swimtime="00:00:00.00" resultid="18722" heatid="19986" lane="1" entrytime="00:03:06.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-06-29" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="347685" swrid="5031429" athleteid="16529">
              <RESULTS>
                <RESULT eventid="3547" points="277" swimtime="00:00:41.49" resultid="18685" heatid="19839" lane="2" entrytime="00:00:42.43" />
                <RESULT eventid="3570" points="179" reactiontime="+91" swimtime="00:03:20.26" resultid="18686" heatid="19876" lane="7" entrytime="00:03:10.05">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="165" swimtime="00:01:42.06" resultid="18687" heatid="19968" lane="3" entrytime="00:01:39.91" />
                <RESULT eventid="3505" points="265" swimtime="00:03:14.27" resultid="18688" heatid="19985" lane="6" entrytime="00:03:09.95">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TWV" nation="AUT" region="TLSV" clubid="15095" swrid="71937" name="Breedy Badger">
          <CONTACT city="Telfs" email="peter.kriegelsteiner@gmx.at" name="Breedy Badger" street="Prof.-A.-Einbergerstraße 28a" zip="6410" />
          <ATHLETES>
            <ATHLETE birthdate="2003-10-30" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41149" swrid="4797185" athleteid="18987">
              <RESULTS>
                <RESULT eventid="3639" points="435" reactiontime="+88" swimtime="00:02:46.42" resultid="18988" heatid="19818" lane="2" entrytime="00:02:46.73">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="489" swimtime="00:00:30.11" resultid="18989" heatid="19934" lane="3" entrytime="00:00:29.75" />
                <RESULT eventid="3555" points="446" reactiontime="+83" swimtime="00:01:13.32" resultid="18990" heatid="19973" lane="7" entrytime="00:01:13.65" />
                <RESULT eventid="3617" points="478" swimtime="00:00:32.06" resultid="18991" heatid="20030" lane="6" entrytime="00:00:31.60" />
                <RESULT eventid="3586" points="380" swimtime="00:02:48.07" resultid="18992" heatid="20064" lane="5" entrytime="00:02:43.37">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="433" reactiontime="+77" swimtime="00:01:08.80" resultid="18993" heatid="20094" lane="6" entrytime="00:01:08.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-09-06" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43493" swrid="5101395" athleteid="19001">
              <RESULTS>
                <RESULT eventid="3547" points="145" swimtime="00:00:51.42" resultid="19002" heatid="19834" lane="3" />
                <RESULT eventid="3621" points="166" swimtime="00:01:57.06" resultid="19003" heatid="19853" lane="4" entrytime="00:01:51.93" />
                <RESULT eventid="3570" points="146" swimtime="00:03:34.43" resultid="19004" heatid="19874" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="210" swimtime="00:00:39.90" resultid="19005" heatid="19921" lane="6" entrytime="00:00:40.91" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-04-19" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="33808" swrid="4075390" athleteid="19047">
              <RESULTS>
                <RESULT eventid="3551" points="578" swimtime="00:00:28.85" resultid="19048" heatid="19852" lane="1" entrytime="00:00:29.36" />
                <RESULT eventid="3649" points="704" reactiontime="+53" swimtime="00:01:54.61" resultid="19049" heatid="19899" lane="4" entrytime="00:01:52.44">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="662" swimtime="00:00:23.99" resultid="19050" heatid="19958" lane="4" entrytime="00:00:23.27" />
                <RESULT eventid="3613" points="658" swimtime="00:00:25.78" resultid="19051" heatid="20039" lane="5" entrytime="00:00:25.69" />
                <RESULT eventid="3530" points="726" reactiontime="+67" swimtime="00:00:52.19" resultid="19052" heatid="20112" lane="4" entrytime="00:00:50.60" />
                <RESULT eventid="15921" points="601" swimtime="00:00:24.77" resultid="20209" heatid="20121" lane="4" late="yes" />
                <RESULT eventid="15972" points="583" swimtime="00:00:25.03" resultid="20210" heatid="20123" lane="4" late="yes" />
                <RESULT eventid="15975" points="553" swimtime="00:00:25.46" resultid="20211" heatid="20125" lane="4" late="yes" />
                <RESULT eventid="15978" points="560" swimtime="00:00:25.36" resultid="20212" heatid="20127" lane="4" late="yes" />
                <RESULT eventid="15981" points="564" swimtime="00:00:25.30" resultid="20213" heatid="20129" lane="4" late="yes" />
                <RESULT eventid="15984" points="531" swimtime="00:00:25.81" resultid="20214" heatid="20131" lane="4" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-08-08" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38126" swrid="4234308" athleteid="19025">
              <RESULTS>
                <RESULT eventid="3639" points="312" reactiontime="+74" swimtime="00:03:05.97" resultid="19026" heatid="19812" lane="4" entrytime="00:03:06.92">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="340" reactiontime="+68" swimtime="00:01:32.30" resultid="19027" heatid="19860" lane="7" entrytime="00:01:28.12" />
                <RESULT eventid="3590" points="361" swimtime="00:00:33.31" resultid="19028" heatid="19928" lane="3" entrytime="00:00:32.84" />
                <RESULT eventid="3555" points="251" reactiontime="+69" swimtime="00:01:28.79" resultid="19029" heatid="19970" lane="6" entrytime="00:01:25.46" />
                <RESULT eventid="3617" points="317" swimtime="00:00:36.74" resultid="19030" heatid="20028" lane="7" entrytime="00:00:35.14" />
                <RESULT eventid="3658" points="305" reactiontime="+74" swimtime="00:05:54.99" resultid="19031" heatid="20042" lane="8" entrytime="00:06:10.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.72" />
                    <SPLIT distance="200" swimtime="00:02:53.43" />
                    <SPLIT distance="300" swimtime="00:04:25.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="388" swimtime="00:00:40.85" resultid="19032" heatid="20073" lane="4" entrytime="00:00:40.05" />
                <RESULT eventid="3636" points="306" swimtime="00:06:39.77" resultid="19033" heatid="20113" lane="3" entrytime="00:06:50.66">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.29" />
                    <SPLIT distance="200" swimtime="00:03:21.28" />
                    <SPLIT distance="300" swimtime="00:05:11.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-05-27" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="33628" swrid="4075350" athleteid="19096">
              <RESULTS>
                <RESULT eventid="3551" points="495" swimtime="00:00:30.38" resultid="19097" heatid="19850" lane="5" entrytime="00:00:31.96" />
                <RESULT eventid="3649" points="559" reactiontime="+73" swimtime="00:02:03.82" resultid="19098" heatid="19899" lane="2" entrytime="00:01:59.79">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="474" reactiontime="+68" swimtime="00:01:03.87" resultid="19099" heatid="19981" lane="4" entrytime="00:01:01.10" />
                <RESULT eventid="3578" points="557" reactiontime="+69" swimtime="00:04:27.32" resultid="19100" heatid="20058" lane="6" entrytime="00:04:17.55">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.83" />
                    <SPLIT distance="200" swimtime="00:02:12.65" />
                    <SPLIT distance="300" swimtime="00:03:19.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="593" reactiontime="+63" swimtime="00:00:55.81" resultid="19101" heatid="20111" lane="4" entrytime="00:00:55.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-29" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="42251" swrid="5082229" athleteid="19068">
              <RESULTS>
                <RESULT eventid="3551" points="137" swimtime="00:00:46.59" resultid="19069" heatid="19848" lane="8" entrytime="00:00:41.61" />
                <RESULT eventid="3594" points="183" swimtime="00:00:36.79" resultid="19070" heatid="19948" lane="2" entrytime="00:00:36.28" />
                <RESULT eventid="3613" points="162" swimtime="00:00:41.12" resultid="19071" heatid="20034" lane="2" entrytime="00:00:40.92" />
                <RESULT eventid="3519" points="160" swimtime="00:00:49.04" resultid="19072" heatid="20079" lane="6" entrytime="00:00:46.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-06-04" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="33999" swrid="4201331" athleteid="19178">
              <RESULTS>
                <RESULT eventid="3590" points="601" swimtime="00:00:28.11" resultid="19179" heatid="19936" lane="3" entrytime="00:00:28.27" />
                <RESULT eventid="3555" points="568" reactiontime="+64" swimtime="00:01:07.66" resultid="19180" heatid="19975" lane="1" entrytime="00:01:08.11" />
                <RESULT eventid="3598" points="445" swimtime="00:01:16.12" resultid="19181" heatid="20010" lane="4" entrytime="00:01:13.80" />
                <RESULT eventid="3617" points="537" swimtime="00:00:30.83" resultid="19182" heatid="20031" lane="2" entrytime="00:00:30.24" />
                <RESULT eventid="3586" points="456" reactiontime="+76" swimtime="00:02:38.21" resultid="19183" heatid="20065" lane="1" entrytime="00:02:41.08">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="530" reactiontime="+78" swimtime="00:01:04.34" resultid="19184" heatid="20099" lane="2" entrytime="00:01:02.65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-12-21" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41842" swrid="4982376" athleteid="19085">
              <RESULTS>
                <RESULT eventid="3551" points="189" swimtime="00:00:41.82" resultid="19086" heatid="19847" lane="1" entrytime="00:00:43.05" />
                <RESULT eventid="3649" points="213" reactiontime="+58" swimtime="00:02:50.73" resultid="19087" heatid="19889" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="208" swimtime="00:00:35.25" resultid="19088" heatid="19949" lane="3" entrytime="00:00:34.93" />
                <RESULT eventid="3613" points="225" swimtime="00:00:36.87" resultid="19089" heatid="20034" lane="8" entrytime="00:00:42.34" />
                <RESULT eventid="3530" points="236" reactiontime="+59" swimtime="00:01:15.87" resultid="19090" heatid="20101" lane="6" entrytime="00:01:21.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-03-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41064" swrid="4925065" athleteid="18057">
              <RESULTS>
                <RESULT eventid="3590" points="242" swimtime="00:00:38.06" resultid="18059" heatid="19923" lane="1" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="3639" points="247" swimtime="00:03:20.86" resultid="19708" heatid="19812" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="258" swimtime="00:02:57.45" resultid="19709" heatid="19878" lane="4" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3505" points="262" swimtime="00:03:14.81" resultid="19710" heatid="19984" lane="6" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="216" swimtime="00:01:36.76" resultid="19711" heatid="20004" lane="1" entrytime="00:01:33.00" />
                <RESULT eventid="3658" points="286" swimtime="00:06:02.57" resultid="19712" heatid="20042" lane="1" entrytime="00:06:09.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.17" />
                    <SPLIT distance="200" swimtime="00:02:57.80" />
                    <SPLIT distance="300" swimtime="00:04:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="252" swimtime="00:01:22.36" resultid="19713" heatid="20087" lane="7" entrytime="00:01:22.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-07-29" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="200183" athleteid="19034">
              <RESULTS>
                <RESULT eventid="3639" points="461" swimtime="00:02:43.22" resultid="19035" heatid="19819" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="488" swimtime="00:00:30.13" resultid="19036" heatid="19935" lane="8" entrytime="00:00:29.60" />
                <RESULT eventid="3555" points="494" reactiontime="+77" swimtime="00:01:10.87" resultid="19037" heatid="19974" lane="7" entrytime="00:01:10.00" />
                <RESULT eventid="3598" points="468" swimtime="00:01:14.83" resultid="19038" heatid="20012" lane="1" entrytime="00:01:11.00" />
                <RESULT eventid="3617" points="496" swimtime="00:00:31.67" resultid="19039" heatid="20030" lane="5" entrytime="00:00:31.40" />
                <RESULT eventid="3523" points="497" reactiontime="+78" swimtime="00:01:05.73" resultid="19040" heatid="20098" lane="1" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-23" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="30137" swrid="4075369" athleteid="19142">
              <RESULTS>
                <RESULT eventid="9711" points="717" reactiontime="+64" swimtime="00:02:07.34" resultid="19143" heatid="19832" lane="5" entrytime="00:02:07.66">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="545" swimtime="00:00:29.43" resultid="19144" heatid="19852" lane="5" entrytime="00:00:27.58" />
                <RESULT eventid="3594" points="614" swimtime="00:00:24.60" resultid="19145" heatid="19957" lane="5" entrytime="00:00:24.34" />
                <RESULT eventid="3605" points="586" swimtime="00:01:02.04" resultid="19146" heatid="20022" lane="5" entrytime="00:00:59.63" />
                <RESULT eventid="1081" points="623" reactiontime="+65" swimtime="00:04:45.38" resultid="19147" heatid="20119" lane="4" entrytime="00:04:41.33">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="200" swimtime="00:02:17.91" />
                    <SPLIT distance="300" swimtime="00:03:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15921" points="592" swimtime="00:00:24.89" resultid="20237" heatid="20121" lane="2" late="yes" />
                <RESULT eventid="15972" points="565" swimtime="00:00:25.29" resultid="20238" heatid="20123" lane="2" late="yes" />
                <RESULT eventid="15975" points="543" swimtime="00:00:25.63" resultid="20239" heatid="20125" lane="2" late="yes" />
                <RESULT eventid="15978" points="512" swimtime="00:00:26.13" resultid="20240" heatid="20127" lane="2" late="yes" />
                <RESULT eventid="15981" points="513" swimtime="00:00:26.11" resultid="20241" heatid="20129" lane="2" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-09-07" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="34029" swrid="4426790" athleteid="18062">
              <RESULTS>
                <RESULT eventid="3590" points="356" swimtime="00:00:33.47" resultid="18063" heatid="19928" lane="8" entrytime="00:00:33.37" entrycourse="LCM" />
                <RESULT eventid="3505" points="350" swimtime="00:02:56.96" resultid="18064" heatid="19989" lane="8" entrytime="00:02:51.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="334" swimtime="00:01:23.74" resultid="18065" heatid="20008" lane="3" entrytime="00:01:20.52" entrycourse="SCM" />
                <RESULT eventid="3658" points="304" swimtime="00:05:55.65" resultid="18066" heatid="20044" lane="5" entrytime="00:05:36.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.32" />
                    <SPLIT distance="200" swimtime="00:02:51.65" />
                    <SPLIT distance="300" swimtime="00:04:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="339" reactiontime="+87" swimtime="00:01:14.66" resultid="18067" heatid="20092" lane="6" entrytime="00:01:10.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-05-23" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="33926" swrid="4790101" athleteid="18953">
              <RESULTS>
                <RESULT eventid="3551" points="595" swimtime="00:00:28.57" resultid="18954" heatid="19852" lane="3" entrytime="00:00:28.13" />
                <RESULT eventid="3649" points="559" reactiontime="+58" swimtime="00:02:03.79" resultid="18955" heatid="19895" lane="5" entrytime="00:02:14.73">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="543" swimtime="00:00:25.62" resultid="18956" heatid="19957" lane="6" entrytime="00:00:25.61" />
                <RESULT eventid="3512" points="410" swimtime="00:02:30.63" resultid="18957" heatid="20000" lane="6" entrytime="00:02:23.06">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="513" swimtime="00:01:04.88" resultid="18958" heatid="20022" lane="3" entrytime="00:01:00.12" />
                <RESULT eventid="3578" points="264" reactiontime="+67" swimtime="00:05:43.05" resultid="18959" heatid="20051" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.35" />
                    <SPLIT distance="200" swimtime="00:02:47.01" />
                    <SPLIT distance="300" swimtime="00:04:20.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" status="DNS" swimtime="00:00:00.00" resultid="18960" heatid="20111" lane="3" entrytime="00:00:55.81" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-12-21" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="44798" athleteid="18936">
              <RESULTS>
                <RESULT eventid="3551" points="337" swimtime="00:00:34.52" resultid="18937" heatid="19845" lane="7" />
                <RESULT eventid="3628" points="335" reactiontime="+71" swimtime="00:01:24.28" resultid="18938" heatid="19864" lane="1" />
                <RESULT eventid="3594" points="411" swimtime="00:00:28.12" resultid="18939" heatid="19946" lane="1" />
                <RESULT eventid="3519" points="391" swimtime="00:00:36.47" resultid="18940" heatid="20076" lane="5" />
                <RESULT eventid="3530" points="322" reactiontime="+71" swimtime="00:01:08.39" resultid="18941" heatid="20100" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-05-14" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="37982" swrid="4329607" athleteid="19073">
              <RESULTS>
                <RESULT eventid="3551" points="294" swimtime="00:00:36.14" resultid="19074" heatid="19845" lane="1" />
                <RESULT eventid="3628" points="345" swimtime="00:01:23.48" resultid="19075" heatid="19868" lane="5" entrytime="00:01:24.36" />
                <RESULT eventid="3594" points="381" swimtime="00:00:28.83" resultid="19076" heatid="19952" lane="3" entrytime="00:00:30.07" />
                <RESULT eventid="3613" points="341" swimtime="00:00:32.08" resultid="19077" heatid="20035" lane="6" entrytime="00:00:33.56" />
                <RESULT eventid="3519" points="386" swimtime="00:00:36.61" resultid="19078" heatid="20082" lane="2" entrytime="00:00:38.33" />
                <RESULT eventid="3530" points="383" reactiontime="+77" swimtime="00:01:04.59" resultid="19079" heatid="20107" lane="6" entrytime="00:01:05.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-02-15" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38536" swrid="4329604" athleteid="19013">
              <RESULTS>
                <RESULT eventid="3639" points="339" reactiontime="+58" swimtime="00:03:00.82" resultid="19014" heatid="19816" lane="1" entrytime="00:02:55.56">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="415" swimtime="00:00:36.27" resultid="19015" heatid="19842" lane="6" entrytime="00:00:35.76" />
                <RESULT eventid="3570" points="328" reactiontime="+59" swimtime="00:02:43.79" resultid="19016" heatid="19882" lane="2" entrytime="00:02:32.72">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" status="DNS" swimtime="00:00:00.00" resultid="19017" heatid="19904" lane="5" />
                <RESULT eventid="3505" status="DNS" swimtime="00:00:00.00" resultid="19018" heatid="19989" lane="7" entrytime="00:02:49.65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-06-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="35110" swrid="4126998" athleteid="19192">
              <RESULTS>
                <RESULT eventid="3639" points="386" reactiontime="+72" swimtime="00:02:53.17" resultid="19193" heatid="19817" lane="1" entrytime="00:02:51.63">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="378" swimtime="00:00:37.41" resultid="19194" heatid="19841" lane="5" entrytime="00:00:36.75" />
                <RESULT eventid="3590" points="424" swimtime="00:00:31.57" resultid="19195" heatid="19933" lane="3" entrytime="00:00:30.10" />
                <RESULT eventid="3598" points="346" swimtime="00:01:22.72" resultid="19196" heatid="20009" lane="8" entrytime="00:01:19.33" />
                <RESULT eventid="3617" points="338" swimtime="00:00:35.97" resultid="19197" heatid="20028" lane="5" entrytime="00:00:34.19" />
                <RESULT eventid="3523" points="387" reactiontime="+77" swimtime="00:01:11.45" resultid="19198" heatid="20096" lane="5" entrytime="00:01:05.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-06-15" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41886" swrid="4600871" athleteid="18994">
              <RESULTS>
                <RESULT eventid="3547" points="201" swimtime="00:00:46.12" resultid="18995" heatid="19838" lane="8" entrytime="00:00:45.15" />
                <RESULT eventid="3570" points="189" swimtime="00:03:16.86" resultid="18996" heatid="19876" lane="2" entrytime="00:03:09.53">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="230" swimtime="00:00:38.72" resultid="18997" heatid="19922" lane="1" entrytime="00:00:40.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-11-02" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="37748" swrid="4909569" athleteid="18049">
              <RESULTS>
                <RESULT eventid="3639" points="437" reactiontime="+85" swimtime="00:02:46.14" resultid="18050" heatid="19820" lane="6" entrytime="00:02:37.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="504" reactiontime="+69" swimtime="00:01:20.94" resultid="18051" heatid="19863" lane="2" entrytime="00:01:18.04" entrycourse="SCM" />
                <RESULT eventid="3538" points="476" reactiontime="+79" swimtime="00:02:59.42" resultid="18052" heatid="19910" lane="7" entrytime="00:02:48.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="388" reactiontime="+76" swimtime="00:01:16.81" resultid="18053" heatid="19974" lane="8" entrytime="00:01:10.95" entrycourse="SCM" />
                <RESULT eventid="3617" points="512" swimtime="00:00:31.32" resultid="18054" heatid="20030" lane="7" entrytime="00:00:31.91" entrycourse="SCM" />
                <RESULT eventid="3514" points="544" swimtime="00:00:36.49" resultid="18055" heatid="20075" lane="6" entrytime="00:00:36.87" entrycourse="SCM" />
                <RESULT eventid="3523" points="436" reactiontime="+75" swimtime="00:01:08.63" resultid="18056" heatid="20097" lane="1" entrytime="00:01:05.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-13" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="24803" swrid="4075532" athleteid="18942">
              <RESULTS>
                <RESULT eventid="3594" points="521" swimtime="00:00:25.97" resultid="18943" heatid="19958" lane="6" entrytime="00:00:25.43" />
                <RESULT eventid="3562" points="445" reactiontime="+74" swimtime="00:01:05.21" resultid="18944" heatid="19980" lane="6" entrytime="00:01:05.01" />
                <RESULT eventid="3613" points="503" swimtime="00:00:28.19" resultid="18945" heatid="20038" lane="5" entrytime="00:00:28.39" />
                <RESULT eventid="3530" points="537" reactiontime="+72" swimtime="00:00:57.71" resultid="18946" heatid="20111" lane="8" entrytime="00:00:57.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-04-13" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41031" swrid="4942827" athleteid="18042">
              <RESULTS>
                <RESULT eventid="3639" points="233" swimtime="00:03:24.89" resultid="18043" heatid="19810" lane="3" entrytime="00:03:22.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="233" swimtime="00:00:43.94" resultid="18044" heatid="19838" lane="6" entrytime="00:00:44.01" entrycourse="SCM" />
                <RESULT eventid="3590" points="248" swimtime="00:00:37.76" resultid="18045" heatid="19923" lane="3" entrytime="00:00:37.26" entrycourse="LCM" />
                <RESULT eventid="3505" points="230" swimtime="00:03:23.58" resultid="18046" heatid="19984" lane="5" entrytime="00:03:15.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="218" swimtime="00:01:36.43" resultid="18047" heatid="20004" lane="5" entrytime="00:01:31.34" entrycourse="SCM" />
                <RESULT eventid="3523" points="199" reactiontime="+72" swimtime="00:01:29.13" resultid="18048" heatid="20087" lane="8" entrytime="00:01:23.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-03-03" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41882" swrid="4992325" athleteid="19119">
              <RESULTS>
                <RESULT eventid="3621" points="313" reactiontime="+80" swimtime="00:01:34.89" resultid="19120" heatid="19855" lane="1" entrytime="00:01:43.33" />
                <RESULT eventid="3555" points="241" reactiontime="+59" swimtime="00:01:30.07" resultid="19121" heatid="19969" lane="3" entrytime="00:01:31.78" />
                <RESULT eventid="3658" points="346" reactiontime="+61" swimtime="00:05:40.60" resultid="19122" heatid="20043" lane="3" entrytime="00:05:53.29">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.60" />
                    <SPLIT distance="200" swimtime="00:02:48.00" />
                    <SPLIT distance="300" swimtime="00:04:15.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="389" swimtime="00:01:11.32" resultid="19123" heatid="20090" lane="3" entrytime="00:01:14.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-10-30" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="42569" swrid="5046056" athleteid="19102">
              <RESULTS>
                <RESULT eventid="3605" points="122" swimtime="00:01:44.58" resultid="19103" heatid="20013" lane="3" entrytime="00:01:41.01" />
                <RESULT eventid="3613" points="60" swimtime="00:00:57.06" resultid="19104" heatid="20032" lane="2" />
                <RESULT eventid="3519" points="139" swimtime="00:00:51.41" resultid="19105" heatid="20077" lane="8" entrytime="00:01:01.37" />
                <RESULT eventid="3530" points="114" reactiontime="+66" swimtime="00:01:36.52" resultid="19106" heatid="20100" lane="6" entrytime="00:01:44.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-09" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38678" swrid="4858660" athleteid="18075">
              <RESULTS>
                <RESULT eventid="3547" points="488" swimtime="00:00:34.37" resultid="18076" heatid="19844" lane="8" entrytime="00:00:33.28" entrycourse="SCM" />
                <RESULT eventid="3570" points="412" swimtime="00:02:31.76" resultid="18077" heatid="19883" lane="4" entrytime="00:02:27.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="426" swimtime="00:00:31.53" resultid="18078" heatid="19932" lane="5" entrytime="00:00:30.54" entrycourse="SCM" />
                <RESULT eventid="3505" points="454" swimtime="00:02:42.29" resultid="18079" heatid="19993" lane="6" entrytime="00:02:29.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="469" swimtime="00:01:14.80" resultid="18080" heatid="20012" lane="2" entrytime="00:01:10.06" entrycourse="SCM" />
                <RESULT eventid="3658" points="387" reactiontime="+65" swimtime="00:05:28.03" resultid="18081" heatid="20046" lane="4" entrytime="00:05:10.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="200" swimtime="00:02:38.22" />
                    <SPLIT distance="300" swimtime="00:04:04.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="402" reactiontime="+75" swimtime="00:01:10.52" resultid="18082" heatid="20095" lane="1" entrytime="00:01:07.74" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-09-07" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41185" swrid="5071972" athleteid="19058">
              <RESULTS>
                <RESULT eventid="3628" points="313" reactiontime="+73" swimtime="00:01:26.21" resultid="19059" heatid="19869" lane="2" entrytime="00:01:23.00" />
                <RESULT eventid="3649" points="314" reactiontime="+81" swimtime="00:02:29.92" resultid="19060" heatid="19893" lane="4" entrytime="00:02:24.93">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3545" points="312" swimtime="00:03:07.56" resultid="19061" heatid="19914" lane="5" entrytime="00:02:57.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="187" swimtime="00:01:27.02" resultid="19062" heatid="19977" lane="4" entrytime="00:01:20.19" />
                <RESULT eventid="3605" points="242" swimtime="00:01:23.34" resultid="19063" heatid="20018" lane="1" entrytime="00:01:17.71" />
                <RESULT eventid="3578" points="353" swimtime="00:05:11.21" resultid="19064" heatid="20055" lane="3" entrytime="00:05:02.54">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.32" />
                    <SPLIT distance="200" swimtime="00:02:33.23" />
                    <SPLIT distance="300" swimtime="00:03:53.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="296" swimtime="00:00:40.00" resultid="19065" heatid="20082" lane="8" entrytime="00:00:38.69" />
                <RESULT eventid="3530" points="322" swimtime="00:01:08.43" resultid="19066" heatid="20106" lane="5" entrytime="00:01:07.27" />
                <RESULT eventid="1081" points="279" swimtime="00:06:12.76" resultid="19067" heatid="20116" lane="4" entrytime="00:06:14.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.17" />
                    <SPLIT distance="200" swimtime="00:03:13.13" />
                    <SPLIT distance="300" swimtime="00:04:53.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-12-05" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38703" swrid="4797183" athleteid="18068">
              <RESULTS>
                <RESULT eventid="3639" points="392" reactiontime="+74" swimtime="00:02:52.23" resultid="18069" heatid="19818" lane="6" entrytime="00:02:46.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="426" swimtime="00:01:25.60" resultid="18070" heatid="19862" lane="4" entrytime="00:01:19.52" entrycourse="SCM" />
                <RESULT eventid="3570" points="385" reactiontime="+74" swimtime="00:02:35.22" resultid="18071" heatid="19874" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="463" swimtime="00:00:30.66" resultid="18072" heatid="19932" lane="2" entrytime="00:00:30.79" entrycourse="LCM" />
                <RESULT eventid="3514" points="490" swimtime="00:00:37.79" resultid="18073" heatid="20074" lane="3" entrytime="00:00:37.41" entrycourse="LCM" />
                <RESULT eventid="3523" points="432" reactiontime="+58" swimtime="00:01:08.84" resultid="18074" heatid="20097" lane="7" entrytime="00:01:05.52" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-24" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="20293" swrid="4102511" athleteid="18998">
              <RESULTS>
                <RESULT eventid="9711" points="370" reactiontime="+85" swimtime="00:02:38.77" resultid="18999" heatid="19829" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="397" reactiontime="+69" swimtime="00:02:18.67" resultid="19000" heatid="19895" lane="1" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-05-18" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="33261" swrid="4075490" athleteid="19185">
              <RESULTS>
                <RESULT eventid="3649" points="591" reactiontime="+50" swimtime="00:02:01.54" resultid="19186" heatid="19899" lane="1" entrytime="00:02:00.40">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="623" swimtime="00:00:24.47" resultid="19187" heatid="19959" lane="5" entrytime="00:00:23.97" />
                <RESULT eventid="3562" points="476" reactiontime="+63" swimtime="00:01:03.78" resultid="19188" heatid="19982" lane="3" entrytime="00:00:57.91" />
                <RESULT eventid="3613" points="611" swimtime="00:00:26.42" resultid="19189" heatid="20039" lane="4" entrytime="00:00:25.41" />
                <RESULT eventid="3519" points="621" swimtime="00:00:31.26" resultid="19190" heatid="20084" lane="6" entrytime="00:00:30.74" />
                <RESULT eventid="3530" points="447" reactiontime="+61" swimtime="00:01:01.35" resultid="19191" heatid="20112" lane="2" entrytime="00:00:53.53" />
                <RESULT eventid="15975" points="521" swimtime="00:00:25.98" resultid="20220" heatid="20125" lane="5" late="yes" />
                <RESULT eventid="15972" points="562" swimtime="00:00:25.33" resultid="20221" heatid="20123" lane="5" late="yes" />
                <RESULT eventid="15921" points="595" swimtime="00:00:24.85" resultid="20222" heatid="20121" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-09" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="35441" swrid="4383150" athleteid="19091">
              <RESULTS>
                <RESULT eventid="3649" points="376" reactiontime="+80" swimtime="00:02:21.20" resultid="19092" heatid="19895" lane="6" entrytime="00:02:16.87">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="442" swimtime="00:00:27.43" resultid="19093" heatid="19957" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="3578" points="365" reactiontime="+78" swimtime="00:05:07.80" resultid="19094" heatid="20055" lane="2" entrytime="00:05:10.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="200" swimtime="00:02:33.31" />
                    <SPLIT distance="300" swimtime="00:03:50.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="437" reactiontime="+77" swimtime="00:01:01.79" resultid="19095" heatid="20109" lane="4" entrytime="00:00:59.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-02-27" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="37221" swrid="4075371" athleteid="19148">
              <RESULTS>
                <RESULT eventid="3590" points="422" swimtime="00:00:31.62" resultid="19149" heatid="19933" lane="7" entrytime="00:00:30.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-10-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41881" swrid="4992324" athleteid="19113">
              <RESULTS>
                <RESULT eventid="3649" points="346" reactiontime="+75" swimtime="00:02:25.16" resultid="19114" heatid="19893" lane="1" entrytime="00:02:35.31" />
                <RESULT eventid="3594" points="420" swimtime="00:00:27.91" resultid="19115" heatid="19952" lane="1" entrytime="00:00:30.98" />
                <RESULT eventid="3613" points="350" swimtime="00:00:31.81" resultid="19116" heatid="20035" lane="8" entrytime="00:00:35.20" />
                <RESULT eventid="3578" points="330" reactiontime="+78" swimtime="00:05:18.22" resultid="19117" heatid="20054" lane="2" entrytime="00:05:34.61">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.50" />
                    <SPLIT distance="200" swimtime="00:02:34.98" />
                    <SPLIT distance="300" swimtime="00:03:58.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="399" reactiontime="+80" swimtime="00:01:03.69" resultid="19118" heatid="20106" lane="6" entrytime="00:01:07.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-07-08" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40818" swrid="4902497" athleteid="18970">
              <RESULTS>
                <RESULT eventid="3639" points="254" swimtime="00:03:19.11" resultid="18971" heatid="19810" lane="2" entrytime="00:03:24.66">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="253" swimtime="00:01:28.56" resultid="18972" heatid="19969" lane="2" entrytime="00:01:32.68" />
                <RESULT eventid="3617" points="309" swimtime="00:00:37.08" resultid="18973" heatid="20026" lane="2" entrytime="00:00:40.69" />
                <RESULT eventid="3658" points="269" reactiontime="+103" swimtime="00:06:10.39" resultid="18974" heatid="20041" lane="5" entrytime="00:06:11.04">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.56" />
                    <SPLIT distance="200" swimtime="00:03:03.36" />
                    <SPLIT distance="300" swimtime="00:04:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="275" swimtime="00:01:20.02" resultid="18975" heatid="20086" lane="5" entrytime="00:01:25.13" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-09-23" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43492" athleteid="20273">
              <RESULTS>
                <RESULT eventid="3617" points="186" swimtime="00:00:43.89" resultid="20274" heatid="20025" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-04-25" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="44185" swrid="5180809" athleteid="19174">
              <RESULTS>
                <RESULT eventid="3547" points="125" swimtime="00:00:54.07" resultid="19175" heatid="19835" lane="2" entrytime="00:00:59.68" />
                <RESULT eventid="3590" points="169" swimtime="00:00:42.92" resultid="19176" heatid="19920" lane="8" entrytime="00:00:46.39" />
                <RESULT eventid="3514" points="148" swimtime="00:00:56.33" resultid="19177" heatid="20069" lane="2" entrytime="00:00:56.07" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-03-09" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40819" swrid="4902498" athleteid="19006">
              <RESULTS>
                <RESULT eventid="3639" points="463" swimtime="00:02:42.99" resultid="19007" heatid="19816" lane="3" entrytime="00:02:52.94">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="396" swimtime="00:00:36.83" resultid="19008" heatid="19841" lane="7" entrytime="00:00:37.52" />
                <RESULT eventid="3570" points="505" swimtime="00:02:21.79" resultid="19009" heatid="19885" lane="5" entrytime="00:02:22.33">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="440" swimtime="00:00:31.18" resultid="19010" heatid="19929" lane="7" entrytime="00:00:32.16" />
                <RESULT eventid="3658" points="487" reactiontime="+72" swimtime="00:05:03.89" resultid="19011" heatid="20048" lane="1" entrytime="00:05:03.67">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="200" swimtime="00:02:28.07" />
                    <SPLIT distance="300" swimtime="00:03:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="454" reactiontime="+48" swimtime="00:01:07.72" resultid="19012" heatid="20094" lane="3" entrytime="00:01:08.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-09-16" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42905" swrid="5087779" athleteid="19137">
              <RESULTS>
                <RESULT eventid="3547" points="141" swimtime="00:00:51.93" resultid="19138" heatid="19835" lane="8" entrytime="00:01:00.16" />
                <RESULT eventid="3590" points="151" swimtime="00:00:44.49" resultid="19139" heatid="19919" lane="8" entrytime="00:00:52.86" />
                <RESULT eventid="3617" points="81" swimtime="00:00:57.94" resultid="19140" heatid="20023" lane="2" />
                <RESULT eventid="3514" points="240" swimtime="00:00:47.92" resultid="19141" heatid="20069" lane="5" entrytime="00:00:54.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-06-28" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="38124" swrid="4736703" athleteid="19124">
              <RESULTS>
                <RESULT eventid="3551" points="198" swimtime="00:00:41.22" resultid="19125" heatid="19846" lane="8" />
                <RESULT eventid="3628" points="301" reactiontime="+60" swimtime="00:01:27.40" resultid="19126" heatid="19867" lane="8" entrytime="00:01:31.33" />
                <RESULT eventid="3545" points="316" reactiontime="+57" swimtime="00:03:06.87" resultid="19127" heatid="19913" lane="8" entrytime="00:03:15.13">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="254" swimtime="00:00:32.99" resultid="19128" heatid="19948" lane="5" entrytime="00:00:35.69" />
                <RESULT eventid="3613" points="204" swimtime="00:00:38.10" resultid="19129" heatid="20032" lane="6" />
                <RESULT eventid="3519" points="304" swimtime="00:00:39.66" resultid="19130" heatid="20080" lane="7" entrytime="00:00:42.97" />
                <RESULT eventid="3530" points="265" swimtime="00:01:13.03" resultid="19131" heatid="20101" lane="4" entrytime="00:01:20.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-27" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="37449" swrid="4487241" athleteid="19053">
              <RESULTS>
                <RESULT eventid="3639" points="476" swimtime="00:02:41.51" resultid="19054" heatid="19819" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="503" reactiontime="+73" swimtime="00:01:21.01" resultid="19055" heatid="19862" lane="2" entrytime="00:01:20.80" />
                <RESULT eventid="3538" points="486" reactiontime="+91" swimtime="00:02:58.19" resultid="19056" heatid="19909" lane="7" entrytime="00:02:57.44">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="403" reactiontime="+90" swimtime="00:01:15.86" resultid="19057" heatid="19972" lane="7" entrytime="00:01:16.93" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-03-27" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40820" swrid="4902499" athleteid="19041">
              <RESULTS>
                <RESULT eventid="3621" points="294" swimtime="00:01:36.89" resultid="19042" heatid="19859" lane="8" entrytime="00:01:31.84" />
                <RESULT eventid="3570" points="337" reactiontime="+73" swimtime="00:02:42.34" resultid="19043" heatid="19879" lane="7" entrytime="00:02:51.29">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="255" swimtime="00:01:28.38" resultid="19044" heatid="19968" lane="4" entrytime="00:01:35.80" />
                <RESULT eventid="3598" points="318" swimtime="00:01:25.07" resultid="19045" heatid="20004" lane="7" entrytime="00:01:32.62" />
                <RESULT eventid="3523" points="390" swimtime="00:01:11.25" resultid="19046" heatid="20087" lane="1" entrytime="00:01:23.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-10-28" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42094" swrid="4982374" athleteid="18036">
              <RESULTS>
                <RESULT eventid="3621" points="408" reactiontime="+67" swimtime="00:01:26.88" resultid="18037" heatid="19861" lane="2" entrytime="00:01:23.44" entrycourse="SCM" />
                <RESULT eventid="3590" points="484" swimtime="00:00:30.22" resultid="18038" heatid="19932" lane="3" entrytime="00:00:30.61" entrycourse="SCM" />
                <RESULT eventid="3617" points="484" swimtime="00:00:31.92" resultid="18039" heatid="20028" lane="3" entrytime="00:00:34.81" entrycourse="LCM" />
                <RESULT eventid="3514" points="437" swimtime="00:00:39.24" resultid="18040" heatid="20073" lane="5" entrytime="00:00:41.05" entrycourse="SCM" />
                <RESULT eventid="3523" points="469" reactiontime="+69" swimtime="00:01:07.00" resultid="18041" heatid="20097" lane="6" entrytime="00:01:05.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-03-27" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40822" swrid="4902500" athleteid="19150">
              <RESULTS>
                <RESULT eventid="3547" points="582" swimtime="00:00:32.40" resultid="19151" heatid="19844" lane="2" entrytime="00:00:32.10" />
                <RESULT eventid="3555" points="531" reactiontime="+63" swimtime="00:01:09.22" resultid="19152" heatid="19974" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="3505" points="496" swimtime="00:02:37.60" resultid="19153" heatid="19993" lane="1" entrytime="00:02:31.62">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="561" swimtime="00:01:10.47" resultid="19154" heatid="20012" lane="7" entrytime="00:01:10.09" />
                <RESULT eventid="3658" points="433" swimtime="00:05:16.01" resultid="19155" heatid="20045" lane="5" entrytime="00:05:24.42">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="200" swimtime="00:02:35.96" />
                    <SPLIT distance="300" swimtime="00:03:57.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3636" points="435" reactiontime="+73" swimtime="00:05:55.35" resultid="19156" heatid="20113" lane="5" entrytime="00:06:36.57">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.29" />
                    <SPLIT distance="200" swimtime="00:02:52.87" />
                    <SPLIT distance="300" swimtime="00:04:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3617" points="587" swimtime="00:00:29.93" resultid="19714" heatid="20031" lane="4" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42629" swrid="5055517" athleteid="18961">
              <RESULTS>
                <RESULT eventid="3514" points="172" swimtime="00:00:53.56" resultid="18962" heatid="20068" lane="4" entrytime="00:00:58.86" />
                <RESULT eventid="3547" points="172" swimtime="00:00:48.65" resultid="18963" heatid="19835" lane="6" entrytime="00:00:59.47" />
                <RESULT eventid="3621" points="160" swimtime="00:01:58.60" resultid="18964" heatid="19853" lane="5" entrytime="00:01:52.60" />
                <RESULT eventid="3570" points="151" swimtime="00:03:32.13" resultid="18965" heatid="19874" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="208" swimtime="00:00:40.04" resultid="18966" heatid="19919" lane="5" entrytime="00:00:47.90" />
                <RESULT eventid="3598" points="170" swimtime="00:01:44.86" resultid="18967" heatid="20002" lane="4" entrytime="00:02:03.53" />
                <RESULT eventid="3617" points="85" swimtime="00:00:56.89" resultid="18968" heatid="20023" lane="7" />
                <RESULT eventid="3523" points="177" reactiontime="+66" swimtime="00:01:32.68" resultid="18969" heatid="20085" lane="4" entrytime="00:01:42.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-10-16" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="44575" swrid="5180808" athleteid="19165">
              <RESULTS>
                <RESULT eventid="3551" points="136" swimtime="00:00:46.67" resultid="19166" heatid="19846" lane="6" entrytime="00:00:46.68" />
                <RESULT eventid="3628" points="264" swimtime="00:01:31.29" resultid="19167" heatid="19865" lane="3" entrytime="00:01:36.62" />
                <RESULT eventid="3649" points="150" reactiontime="+64" swimtime="00:03:11.66" resultid="19168" heatid="19889" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="217" swimtime="00:00:34.76" resultid="19169" heatid="19947" lane="6" entrytime="00:00:39.10" />
                <RESULT eventid="3605" points="134" swimtime="00:01:41.48" resultid="19170" heatid="20013" lane="4" entrytime="00:01:36.89" />
                <RESULT eventid="3613" points="110" swimtime="00:00:46.73" resultid="19171" heatid="20032" lane="7" />
                <RESULT eventid="3519" points="272" swimtime="00:00:41.16" resultid="19172" heatid="20079" lane="5" entrytime="00:00:44.81" />
                <RESULT eventid="3530" points="196" reactiontime="+63" swimtime="00:01:20.72" resultid="19173" heatid="20101" lane="1" entrytime="00:01:25.73" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-02-24" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="40823" swrid="4902501" athleteid="19157">
              <RESULTS>
                <RESULT eventid="3547" points="474" swimtime="00:00:34.69" resultid="19158" heatid="19842" lane="2" entrytime="00:00:35.84" />
                <RESULT eventid="3570" points="393" reactiontime="+66" swimtime="00:02:34.17" resultid="19159" heatid="19879" lane="1" entrytime="00:02:51.91">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="448" swimtime="00:00:31.00" resultid="19160" heatid="19932" lane="7" entrytime="00:00:30.80" />
                <RESULT eventid="3505" points="379" swimtime="00:02:52.32" resultid="19161" heatid="19988" lane="4" entrytime="00:02:51.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="397" swimtime="00:01:19.02" resultid="19162" heatid="20010" lane="1" entrytime="00:01:16.85" />
                <RESULT eventid="3617" points="342" swimtime="00:00:35.84" resultid="19163" heatid="20027" lane="1" entrytime="00:00:37.65" />
                <RESULT eventid="3523" points="396" reactiontime="+63" swimtime="00:01:10.87" resultid="19164" heatid="20095" lane="3" entrytime="00:01:07.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2006-06-21" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="42568" swrid="5046055" athleteid="19080">
              <RESULTS>
                <RESULT eventid="3547" points="197" swimtime="00:00:46.45" resultid="19081" heatid="19836" lane="8" entrytime="00:00:54.23" />
                <RESULT eventid="3590" points="220" swimtime="00:00:39.28" resultid="19082" heatid="19920" lane="6" entrytime="00:00:44.93" />
                <RESULT eventid="3617" points="151" swimtime="00:00:47.03" resultid="19083" heatid="20025" lane="1" entrytime="00:00:44.71" />
                <RESULT eventid="3514" points="200" swimtime="00:00:50.90" resultid="19084" heatid="20069" lane="6" entrytime="00:00:55.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="24804" swrid="4064851" athleteid="18947">
              <RESULTS>
                <RESULT eventid="3649" points="548" reactiontime="+73" swimtime="00:02:04.59" resultid="18948" heatid="19899" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="576" swimtime="00:00:25.13" resultid="18949" heatid="19959" lane="3" entrytime="00:00:24.63" />
                <RESULT eventid="3562" points="540" reactiontime="+75" swimtime="00:01:01.16" resultid="18950" heatid="19982" lane="6" entrytime="00:00:58.17" />
                <RESULT eventid="3613" points="596" swimtime="00:00:26.65" resultid="18951" heatid="20039" lane="6" entrytime="00:00:26.89" />
                <RESULT eventid="3530" points="555" reactiontime="+73" swimtime="00:00:57.05" resultid="18952" heatid="20112" lane="1" entrytime="00:00:54.67" />
                <RESULT eventid="15972" points="496" swimtime="00:00:26.40" resultid="20263" heatid="20123" lane="8" late="yes" />
                <RESULT eventid="15921" points="585" swimtime="00:00:24.99" resultid="20264" heatid="20121" lane="8" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-04-14" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="35371" swrid="4805871" athleteid="19107">
              <RESULTS>
                <RESULT eventid="3551" points="326" swimtime="00:00:34.90" resultid="19108" heatid="19845" lane="2" />
                <RESULT eventid="3649" points="395" reactiontime="+62" swimtime="00:02:18.98" resultid="19109" heatid="19894" lane="7" entrytime="00:02:21.24">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="426" swimtime="00:00:27.78" resultid="19110" heatid="19946" lane="7" />
                <RESULT eventid="3578" points="216" reactiontime="+60" swimtime="00:06:06.31" resultid="19111" heatid="20051" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                    <SPLIT distance="200" swimtime="00:02:48.38" />
                    <SPLIT distance="300" swimtime="00:04:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="455" reactiontime="+63" swimtime="00:01:00.95" resultid="19112" heatid="20109" lane="6" entrytime="00:00:59.86" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-07-28" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="37223" swrid="4287196" athleteid="18981">
              <RESULTS>
                <RESULT eventid="9711" points="428" reactiontime="+72" swimtime="00:02:31.22" resultid="18982" heatid="19832" lane="8" entrytime="00:02:21.06">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="463" reactiontime="+61" swimtime="00:01:15.67" resultid="18983" heatid="19872" lane="1" entrytime="00:01:11.26" />
                <RESULT eventid="3545" points="456" reactiontime="+72" swimtime="00:02:45.31" resultid="18984" heatid="19916" lane="7" entrytime="00:02:35.26">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3578" points="333" reactiontime="+57" swimtime="00:05:17.32" resultid="18985" heatid="20055" lane="4" entrytime="00:04:54.16">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.32" />
                    <SPLIT distance="200" swimtime="00:02:31.61" />
                    <SPLIT distance="300" swimtime="00:03:53.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="515" swimtime="00:00:33.26" resultid="18986" heatid="20084" lane="7" entrytime="00:00:32.87" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-17" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="25995" swrid="4075327" athleteid="19132">
              <RESULTS>
                <RESULT eventid="9711" points="721" reactiontime="+67" swimtime="00:02:07.10" resultid="19133" heatid="19832" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="622" swimtime="00:00:24.49" resultid="19134" heatid="19959" lane="4" entrytime="00:00:23.25" />
                <RESULT eventid="3613" points="638" swimtime="00:00:26.05" resultid="19135" heatid="20039" lane="2" entrytime="00:00:26.95" />
                <RESULT eventid="3530" points="725" reactiontime="+55" swimtime="00:00:52.21" resultid="19136" heatid="20112" lane="5" entrytime="00:00:51.05" />
                <RESULT eventid="15921" points="592" swimtime="00:00:24.90" resultid="20223" heatid="20121" lane="3" late="yes" />
                <RESULT eventid="15972" points="585" swimtime="00:00:25.00" resultid="20224" heatid="20123" lane="3" late="yes" />
                <RESULT eventid="15975" points="558" swimtime="00:00:25.39" resultid="20225" heatid="20125" lane="3" late="yes" />
                <RESULT eventid="15978" points="544" swimtime="00:00:25.61" resultid="20226" heatid="20127" lane="3" late="yes" />
                <RESULT eventid="15981" points="546" swimtime="00:00:25.58" resultid="20227" heatid="20129" lane="3" late="yes" />
                <RESULT eventid="15984" points="569" swimtime="00:00:25.22" resultid="20228" heatid="20131" lane="3" late="yes" />
                <RESULT eventid="15987" points="627" swimtime="00:00:24.43" resultid="20229" heatid="20133" lane="3" late="yes" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="12864" points="656" reactiontime="+62" swimtime="00:03:36.59" resultid="19199" heatid="20137" lane="4" entrytime="00:03:25.08">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.10" />
                    <SPLIT distance="200" swimtime="00:01:47.12" />
                    <SPLIT distance="300" swimtime="00:02:42.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19142" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="19185" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="19132" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="19047" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12820" points="568" swimtime="00:04:10.16" resultid="19201" heatid="20141" lane="4" entrytime="00:03:49.35">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="200" swimtime="00:02:20.19" />
                    <SPLIT distance="300" swimtime="00:03:18.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18953" number="1" />
                    <RELAYPOSITION athleteid="19185" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="19142" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="19047" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="12820" points="533" swimtime="00:04:15.54" resultid="19200" heatid="20140" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="200" swimtime="00:02:19.26" />
                    <SPLIT distance="300" swimtime="00:03:19.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19096" number="1" />
                    <RELAYPOSITION athleteid="18981" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="18947" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="18942" number="4" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="12864" points="577" reactiontime="+61" swimtime="00:03:46.09" resultid="19615" heatid="20136" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.52" />
                    <SPLIT distance="200" swimtime="00:01:51.32" />
                    <SPLIT distance="300" swimtime="00:02:49.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18947" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="18942" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="18953" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="19096" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="12862" points="512" reactiontime="+77" swimtime="00:04:24.51" resultid="19202" heatid="20135" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="200" swimtime="00:02:11.60" />
                    <SPLIT distance="300" swimtime="00:03:18.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19034" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="18036" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="19006" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="19178" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="3574" points="511" swimtime="00:04:50.31" resultid="19204" heatid="20139" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="200" swimtime="00:02:34.79" />
                    <SPLIT distance="300" swimtime="00:03:45.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18075" number="1" />
                    <RELAYPOSITION athleteid="18049" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="19178" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="19034" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="12862" points="429" reactiontime="+74" swimtime="00:04:40.61" resultid="19203" heatid="20134" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="200" swimtime="00:02:19.56" />
                    <SPLIT distance="300" swimtime="00:03:28.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19157" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="18075" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="18049" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="19192" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="3574" points="491" swimtime="00:04:54.20" resultid="19205" heatid="20138" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                    <SPLIT distance="200" swimtime="00:02:36.52" />
                    <SPLIT distance="300" swimtime="00:03:49.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19150" number="1" />
                    <RELAYPOSITION athleteid="18068" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="18987" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="18036" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TSD" nation="AUT" region="VLSV" clubid="13549" swrid="65825" name="Breedy Badger">
          <CONTACT city="Dornbirn" email="Stefanie.Kernbeiss@gmail.com" name="Breedy Badger" state="VB" street="Sebastianstraße 2" zip="6850" />
          <ATHLETES>
            <ATHLETE birthdate="1998-05-19" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="34775" swrid="4254411" athleteid="17224">
              <RESULTS>
                <RESULT eventid="9711" points="391" reactiontime="+69" swimtime="00:02:35.88" resultid="17225" heatid="19828" lane="6" entrytime="00:02:38.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="444" reactiontime="+70" swimtime="00:02:13.69" resultid="17226" heatid="19897" lane="2" entrytime="00:02:08.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="405" swimtime="00:00:28.24" resultid="17227" heatid="19955" lane="2" entrytime="00:00:27.59" entrycourse="LCM" />
                <RESULT eventid="3512" points="385" swimtime="00:02:33.77" resultid="17228" heatid="19999" lane="4" entrytime="00:02:32.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="364" swimtime="00:01:12.71" resultid="17229" heatid="20020" lane="1" entrytime="00:01:11.42" entrycourse="LCM" />
                <RESULT eventid="3578" points="479" swimtime="00:04:41.24" resultid="17230" heatid="20057" lane="4" entrytime="00:04:28.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="200" swimtime="00:02:20.04" />
                    <SPLIT distance="300" swimtime="00:03:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="266" swimtime="00:00:41.44" resultid="17231" heatid="20081" lane="1" entrytime="00:00:40.56" entrycourse="LCM" />
                <RESULT eventid="3530" points="424" reactiontime="+70" swimtime="00:01:02.41" resultid="17232" heatid="20110" lane="7" entrytime="00:00:58.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-11-03" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="34934" swrid="4341719" athleteid="17095">
              <RESULTS>
                <RESULT eventid="3551" points="482" swimtime="00:00:30.65" resultid="17096" heatid="19851" lane="8" entrytime="00:00:31.52" entrycourse="LCM" />
                <RESULT eventid="3649" points="546" reactiontime="+63" swimtime="00:02:04.77" resultid="17097" heatid="19898" lane="1" entrytime="00:02:06.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="476" swimtime="00:00:26.77" resultid="17098" heatid="19956" lane="3" entrytime="00:00:26.98" entrycourse="LCM" />
                <RESULT eventid="3562" points="531" reactiontime="+82" swimtime="00:01:01.49" resultid="17099" heatid="19981" lane="3" entrytime="00:01:02.33" entrycourse="LCM" />
                <RESULT eventid="3605" points="493" swimtime="00:01:05.71" resultid="17100" heatid="20021" lane="3" entrytime="00:01:05.30" entrycourse="LCM" />
                <RESULT eventid="3578" points="561" reactiontime="+76" swimtime="00:04:26.77" resultid="17101" heatid="20058" lane="1" entrytime="00:04:24.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.95" />
                    <SPLIT distance="200" swimtime="00:02:11.18" />
                    <SPLIT distance="300" swimtime="00:03:19.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3588" points="531" reactiontime="+64" swimtime="00:02:17.65" resultid="17102" heatid="20067" lane="5" entrytime="00:02:18.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="526" reactiontime="+82" swimtime="00:05:02.00" resultid="17103" heatid="20119" lane="1" entrytime="00:05:05.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.93" />
                    <SPLIT distance="200" swimtime="00:02:27.10" />
                    <SPLIT distance="300" swimtime="00:03:53.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-03-29" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="38426" swrid="4746943" athleteid="17205">
              <RESULTS>
                <RESULT eventid="9711" points="470" reactiontime="+56" swimtime="00:02:26.60" resultid="17206" heatid="19830" lane="4" entrytime="00:02:28.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3551" points="426" swimtime="00:00:31.94" resultid="17207" heatid="19850" lane="1" entrytime="00:00:32.66" entrycourse="LCM" />
                <RESULT eventid="3545" points="375" reactiontime="+64" swimtime="00:02:56.49" resultid="17208" heatid="19914" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="441" swimtime="00:00:27.47" resultid="17209" heatid="19954" lane="5" entrytime="00:00:27.92" entrycourse="LCM" />
                <RESULT eventid="3512" points="465" swimtime="00:02:24.44" resultid="17210" heatid="20000" lane="1" entrytime="00:02:27.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="477" swimtime="00:01:06.43" resultid="17211" heatid="20021" lane="1" entrytime="00:01:07.12" entrycourse="LCM" />
                <RESULT eventid="3613" points="423" swimtime="00:00:29.87" resultid="17212" heatid="20036" lane="3" entrytime="00:00:31.55" entrycourse="LCM" />
                <RESULT eventid="3530" points="499" reactiontime="+66" swimtime="00:00:59.11" resultid="17213" heatid="20108" lane="6" entrytime="00:01:02.59" entrycourse="LCM" />
                <RESULT eventid="1081" points="487" reactiontime="+71" swimtime="00:05:09.83" resultid="17214" heatid="20118" lane="6" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="200" swimtime="00:02:28.85" />
                    <SPLIT distance="300" swimtime="00:04:02.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-10-25" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38444" swrid="4746938" athleteid="17169">
              <RESULTS>
                <RESULT eventid="3639" points="380" swimtime="00:02:54.09" resultid="17170" heatid="19811" lane="5" entrytime="00:03:15.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="418" reactiontime="+61" swimtime="00:01:26.13" resultid="17171" heatid="19857" lane="6" entrytime="00:01:36.10" entrycourse="LCM" />
                <RESULT eventid="3538" points="412" reactiontime="+74" swimtime="00:03:08.19" resultid="17172" heatid="19905" lane="4" entrytime="00:03:31.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="310" swimtime="00:01:22.77" resultid="17173" heatid="19969" lane="5" entrytime="00:01:30.00" />
                <RESULT eventid="3617" points="335" swimtime="00:00:36.08" resultid="17174" heatid="20026" lane="4" entrytime="00:00:39.87" entrycourse="LCM" />
                <RESULT eventid="3658" points="368" swimtime="00:05:33.63" resultid="17175" heatid="20043" lane="8" entrytime="00:05:57.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="200" swimtime="00:02:42.93" />
                    <SPLIT distance="300" swimtime="00:04:09.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="424" swimtime="00:00:39.65" resultid="17176" heatid="20072" lane="5" entrytime="00:00:43.05" entrycourse="LCM" />
                <RESULT eventid="3523" points="358" reactiontime="+62" swimtime="00:01:13.30" resultid="17177" heatid="20088" lane="6" entrytime="00:01:17.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-07-08" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41365" swrid="4942232" athleteid="17151">
              <RESULTS>
                <RESULT eventid="9711" points="313" reactiontime="+62" swimtime="00:02:47.83" resultid="17152" heatid="19826" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3628" points="290" swimtime="00:01:28.49" resultid="17153" heatid="19866" lane="5" entrytime="00:01:33.33" entrycourse="LCM" />
                <RESULT eventid="3545" points="292" reactiontime="+73" swimtime="00:03:11.68" resultid="17154" heatid="19912" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3512" points="276" swimtime="00:02:51.74" resultid="17155" heatid="19995" lane="6" entrytime="00:03:13.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="293" swimtime="00:01:18.14" resultid="17156" heatid="20014" lane="3" entrytime="00:01:30.29" entrycourse="LCM" />
                <RESULT eventid="3578" points="334" swimtime="00:05:17.06" resultid="17157" heatid="20053" lane="5" entrytime="00:05:49.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="200" swimtime="00:02:34.72" />
                    <SPLIT distance="300" swimtime="00:03:57.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="299" swimtime="00:00:39.84" resultid="17158" heatid="20080" lane="1" entrytime="00:00:43.15" entrycourse="LCM" />
                <RESULT eventid="3530" points="330" reactiontime="+78" swimtime="00:01:07.84" resultid="17159" heatid="20104" lane="7" entrytime="00:01:14.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-05-16" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38056" swrid="4746941" athleteid="17196">
              <RESULTS>
                <RESULT eventid="3639" points="317" reactiontime="+81" swimtime="00:03:04.97" resultid="17197" heatid="19811" lane="7" entrytime="00:03:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="308" swimtime="00:01:35.43" resultid="17198" heatid="19856" lane="4" entrytime="00:01:38.22" entrycourse="LCM" />
                <RESULT eventid="3538" points="302" reactiontime="+80" swimtime="00:03:28.83" resultid="17199" heatid="19906" lane="8" entrytime="00:03:31.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="343" swimtime="00:00:33.87" resultid="17200" heatid="19925" lane="2" entrytime="00:00:35.10" entrycourse="LCM" />
                <RESULT eventid="3598" points="313" swimtime="00:01:25.52" resultid="17201" heatid="20003" lane="5" entrytime="00:01:34.24" entrycourse="LCM" />
                <RESULT eventid="3658" points="313" reactiontime="+75" swimtime="00:05:52.15" resultid="17202" heatid="20043" lane="7" entrytime="00:05:56.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                    <SPLIT distance="200" swimtime="00:02:52.76" />
                    <SPLIT distance="300" swimtime="00:04:25.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="344" swimtime="00:00:42.53" resultid="17203" heatid="20071" lane="5" entrytime="00:00:44.96" entrycourse="LCM" />
                <RESULT eventid="3523" points="321" reactiontime="+70" swimtime="00:01:16.01" resultid="17204" heatid="20088" lane="1" entrytime="00:01:18.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-02-10" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="28946" swrid="4075533" athleteid="17113">
              <RESULTS>
                <RESULT eventid="3519" points="534" swimtime="00:00:32.86" resultid="17114" heatid="20084" lane="2" entrytime="00:00:31.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-08-28" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="34941" swrid="4395263" athleteid="17133">
              <RESULTS>
                <RESULT eventid="3639" points="417" reactiontime="+81" swimtime="00:02:48.74" resultid="17134" heatid="19818" lane="8" entrytime="00:02:48.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="482" reactiontime="+66" swimtime="00:02:24.02" resultid="17135" heatid="19886" lane="1" entrytime="00:02:21.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-10-06" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38427" swrid="4705053" athleteid="17124">
              <RESULTS>
                <RESULT eventid="3639" points="415" swimtime="00:02:49.02" resultid="17125" heatid="19815" lane="3" entrytime="00:02:57.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="428" swimtime="00:01:25.47" resultid="17126" heatid="19858" lane="5" entrytime="00:01:32.35" entrycourse="LCM" />
                <RESULT eventid="3538" points="462" reactiontime="+75" swimtime="00:03:01.13" resultid="17127" heatid="19908" lane="8" entrytime="00:03:11.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="421" swimtime="00:00:31.66" resultid="17128" heatid="19930" lane="6" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="3617" points="351" swimtime="00:00:35.52" resultid="17129" heatid="20027" lane="2" entrytime="00:00:37.45" entrycourse="LCM" />
                <RESULT eventid="3658" points="435" reactiontime="+66" swimtime="00:05:15.51" resultid="17130" heatid="20047" lane="1" entrytime="00:05:10.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="200" swimtime="00:02:38.98" />
                    <SPLIT distance="300" swimtime="00:03:59.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="421" swimtime="00:00:39.76" resultid="17131" heatid="20073" lane="3" entrytime="00:00:41.26" entrycourse="LCM" />
                <RESULT eventid="3523" points="398" swimtime="00:01:10.78" resultid="17132" heatid="20093" lane="3" entrytime="00:01:08.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-09-25" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="38366" swrid="4520479" athleteid="17115">
              <RESULTS>
                <RESULT eventid="9711" points="345" swimtime="00:02:42.46" resultid="17116" heatid="19827" lane="3" entrytime="00:02:49.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="358" reactiontime="+71" swimtime="00:02:23.63" resultid="17117" heatid="19895" lane="8" entrytime="00:02:18.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="354" swimtime="00:00:29.54" resultid="17118" heatid="19952" lane="6" entrytime="00:00:30.11" entrycourse="LCM" />
                <RESULT eventid="3512" points="348" swimtime="00:02:39.09" resultid="17119" heatid="19998" lane="4" entrytime="00:02:38.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="317" swimtime="00:01:16.11" resultid="17120" heatid="20019" lane="1" entrytime="00:01:14.38" entrycourse="LCM" />
                <RESULT eventid="3578" points="396" reactiontime="+70" swimtime="00:04:59.59" resultid="17121" heatid="20056" lane="1" entrytime="00:04:50.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="200" swimtime="00:02:25.48" />
                    <SPLIT distance="300" swimtime="00:03:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3519" points="303" swimtime="00:00:39.69" resultid="17122" heatid="20080" lane="2" entrytime="00:00:42.94" entrycourse="LCM" />
                <RESULT eventid="3530" points="388" reactiontime="+69" swimtime="00:01:04.31" resultid="17123" heatid="20107" lane="4" entrytime="00:01:04.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-17" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="34943" swrid="4395266" athleteid="17178">
              <RESULTS>
                <RESULT eventid="3621" points="474" reactiontime="+63" swimtime="00:01:22.65" resultid="17179" heatid="19863" lane="1" entrytime="00:01:18.56" entrycourse="LCM" />
                <RESULT eventid="3570" points="596" reactiontime="+59" swimtime="00:02:14.24" resultid="17180" heatid="19887" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3538" points="475" reactiontime="+62" swimtime="00:02:59.49" resultid="17181" heatid="19910" lane="2" entrytime="00:02:48.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="524" swimtime="00:00:29.43" resultid="17182" heatid="19935" lane="1" entrytime="00:00:29.26" entrycourse="LCM" />
                <RESULT eventid="3617" points="428" swimtime="00:00:33.25" resultid="17183" heatid="20028" lane="4" entrytime="00:00:34.11" entrycourse="LCM" />
                <RESULT eventid="3658" points="559" reactiontime="+72" swimtime="00:04:50.19" resultid="17184" heatid="20050" lane="1" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="200" swimtime="00:02:20.29" />
                    <SPLIT distance="300" swimtime="00:03:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="498" swimtime="00:00:37.58" resultid="17185" heatid="20075" lane="2" entrytime="00:00:36.90" entrycourse="LCM" />
                <RESULT eventid="3523" points="600" reactiontime="+61" swimtime="00:01:01.71" resultid="17186" heatid="20099" lane="3" entrytime="00:01:01.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-08-21" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="35393" swrid="4364370" athleteid="17142">
              <RESULTS>
                <RESULT eventid="3639" points="504" reactiontime="+75" swimtime="00:02:38.45" resultid="17143" heatid="19820" lane="3" entrytime="00:02:37.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="474" reactiontime="+82" swimtime="00:01:22.66" resultid="17144" heatid="19862" lane="7" entrytime="00:01:20.88" entrycourse="LCM" />
                <RESULT eventid="3538" points="484" reactiontime="+69" swimtime="00:02:58.35" resultid="17145" heatid="19909" lane="4" entrytime="00:02:52.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="412" swimtime="00:01:15.31" resultid="17146" heatid="19972" lane="4" entrytime="00:01:15.70" entrycourse="LCM" />
                <RESULT eventid="3617" points="445" swimtime="00:00:32.82" resultid="17147" heatid="20029" lane="7" entrytime="00:00:33.36" entrycourse="LCM" />
                <RESULT eventid="3658" points="477" reactiontime="+84" swimtime="00:05:06.04" resultid="17148" heatid="20049" lane="1" entrytime="00:04:58.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.52" />
                    <SPLIT distance="200" swimtime="00:02:28.60" />
                    <SPLIT distance="300" swimtime="00:03:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="461" swimtime="00:00:38.56" resultid="17149" heatid="20074" lane="5" entrytime="00:00:37.31" entrycourse="LCM" />
                <RESULT eventid="3523" points="472" reactiontime="+68" swimtime="00:01:06.85" resultid="17150" heatid="20097" lane="2" entrytime="00:01:05.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-04-27" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="AUT" license="41677" swrid="4520495" athleteid="17187">
              <RESULTS>
                <RESULT eventid="3551" points="304" swimtime="00:00:35.74" resultid="17188" heatid="19849" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="3649" points="382" swimtime="00:02:20.56" resultid="17189" heatid="19892" lane="6" entrytime="00:02:40.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="368" swimtime="00:00:29.17" resultid="17190" heatid="19951" lane="6" entrytime="00:00:31.22" entrycourse="LCM" />
                <RESULT eventid="3562" points="352" reactiontime="+81" swimtime="00:01:10.54" resultid="17191" heatid="19977" lane="5" entrytime="00:01:21.41" entrycourse="LCM" />
                <RESULT eventid="3613" points="388" swimtime="00:00:30.74" resultid="17192" heatid="20035" lane="3" entrytime="00:00:33.46" entrycourse="LCM" />
                <RESULT eventid="3578" points="368" reactiontime="+70" swimtime="00:05:06.86" resultid="17193" heatid="20052" lane="3" entrytime="00:06:00.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.82" />
                    <SPLIT distance="200" swimtime="00:02:30.56" />
                    <SPLIT distance="300" swimtime="00:03:49.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3588" points="311" reactiontime="+78" swimtime="00:02:44.43" resultid="17194" heatid="20066" lane="2" entrytime="00:02:53.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3530" points="376" reactiontime="+79" swimtime="00:01:04.96" resultid="17195" heatid="20104" lane="5" entrytime="00:01:13.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-12-29" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="37956" swrid="4520474" athleteid="17104">
              <RESULTS>
                <RESULT eventid="3639" points="420" reactiontime="+67" swimtime="00:02:48.39" resultid="17105" heatid="19815" lane="7" entrytime="00:02:58.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="414" reactiontime="+95" swimtime="00:02:31.58" resultid="17106" heatid="19882" lane="7" entrytime="00:02:32.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="412" swimtime="00:00:31.87" resultid="17107" heatid="19929" lane="8" entrytime="00:00:32.75" entrycourse="LCM" />
                <RESULT eventid="3505" points="376" swimtime="00:02:52.83" resultid="17108" heatid="19987" lane="5" entrytime="00:02:57.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3598" points="377" swimtime="00:01:20.39" resultid="17109" heatid="20007" lane="4" entrytime="00:01:23.28" entrycourse="LCM" />
                <RESULT eventid="3658" points="452" reactiontime="+85" swimtime="00:05:11.52" resultid="17110" heatid="20046" lane="1" entrytime="00:05:16.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.40" />
                    <SPLIT distance="200" swimtime="00:02:34.90" />
                    <SPLIT distance="300" swimtime="00:03:54.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3514" points="338" swimtime="00:00:42.78" resultid="17111" heatid="20072" lane="4" entrytime="00:00:42.80" entrycourse="LCM" />
                <RESULT eventid="3523" points="391" swimtime="00:01:11.16" resultid="17112" heatid="20092" lane="3" entrytime="00:01:10.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-02-24" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="38054" swrid="4520492" athleteid="17160">
              <RESULTS>
                <RESULT eventid="3639" points="360" swimtime="00:02:57.27" resultid="17161" heatid="19816" lane="5" entrytime="00:02:52.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="360" swimtime="00:01:30.58" resultid="17162" heatid="19859" lane="3" entrytime="00:01:29.63" entrycourse="LCM" />
                <RESULT eventid="3538" points="405" reactiontime="+66" swimtime="00:03:09.27" resultid="17163" heatid="19908" lane="1" entrytime="00:03:10.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3555" points="329" swimtime="00:01:21.20" resultid="17164" heatid="19971" lane="2" entrytime="00:01:20.51" entrycourse="LCM" />
                <RESULT eventid="3617" points="334" swimtime="00:00:36.11" resultid="17165" heatid="20028" lane="8" entrytime="00:00:35.93" entrycourse="LCM" />
                <RESULT eventid="3658" points="410" reactiontime="+78" swimtime="00:05:21.69" resultid="17166" heatid="20044" lane="4" entrytime="00:05:35.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="200" swimtime="00:02:38.33" />
                    <SPLIT distance="300" swimtime="00:04:01.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3586" points="274" reactiontime="+66" swimtime="00:03:07.35" resultid="17167" heatid="20063" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3523" points="365" swimtime="00:01:12.86" resultid="17168" heatid="20092" lane="4" entrytime="00:01:10.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="12862" points="421" reactiontime="+82" swimtime="00:04:42.32" resultid="17233" heatid="20135" lane="6" entrytime="00:04:21.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.11" />
                    <SPLIT distance="200" swimtime="00:02:23.41" />
                    <SPLIT distance="300" swimtime="00:03:33.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17124" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="17169" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="17160" number="3" reactiontime="+2" />
                    <RELAYPOSITION athleteid="17104" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="3574" points="449" swimtime="00:05:03.20" resultid="17234" heatid="20139" lane="1" entrytime="00:04:56.21">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.23" />
                    <SPLIT distance="200" swimtime="00:02:44.18" />
                    <SPLIT distance="300" swimtime="00:04:00.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17104" number="1" />
                    <RELAYPOSITION athleteid="17142" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="17133" number="3" />
                    <RELAYPOSITION athleteid="17178" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Julia" gender="F" lastname="Janke-Frosch" license="27440" type="HEADCOACH">
              <CONTACT city="Dornbirn" email="Stefanie.Kernbeiss@gmail.com" state="VB" street="Sebastianstraße 2" zip="6850" />
            </COACH>
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="ROSENH" nation="GER" region="02" clubid="19716" swrid="66109" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="257560" swrid="4406859" athleteid="19717">
              <RESULTS>
                <RESULT eventid="9711" points="343" reactiontime="+71" swimtime="00:02:42.70" resultid="19718" heatid="19830" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3649" points="392" reactiontime="+75" swimtime="00:02:19.30" resultid="19719" heatid="19897" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="352" reactiontime="+61" swimtime="00:01:10.52" resultid="19720" heatid="19981" lane="1" entrytime="00:01:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="372780" swrid="5166325" athleteid="19726">
              <RESULTS>
                <RESULT eventid="3639" points="566" swimtime="00:02:32.44" resultid="19727" heatid="19821" lane="5" entrytime="00:02:34.70">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3547" points="475" swimtime="00:00:34.68" resultid="19728" heatid="19844" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="3570" points="598" reactiontime="+64" swimtime="00:02:14.06" resultid="19729" heatid="19887" lane="2" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="573" swimtime="00:00:28.57" resultid="19730" heatid="19937" lane="2" entrytime="00:00:28.70" />
                <RESULT eventid="3555" points="583" reactiontime="+64" swimtime="00:01:07.07" resultid="19731" heatid="19975" lane="2" entrytime="00:01:07.40" />
                <RESULT eventid="20145" points="578" swimtime="00:00:28.48" resultid="20150" heatid="20148" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="288564" swrid="4155795" athleteid="19765">
              <RESULTS>
                <RESULT eventid="3551" points="414" swimtime="00:00:32.25" resultid="19766" heatid="19851" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="3649" points="374" reactiontime="+72" swimtime="00:02:21.56" resultid="19767" heatid="19897" lane="7" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="459" swimtime="00:00:27.09" resultid="19768" heatid="19957" lane="7" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="200640" swrid="4154598" athleteid="19721">
              <RESULTS>
                <RESULT eventid="3639" points="453" reactiontime="+70" swimtime="00:02:44.23" resultid="19722" heatid="19820" lane="2" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3570" points="481" reactiontime="+71" swimtime="00:02:24.15" resultid="19723" heatid="19887" lane="8" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="559" swimtime="00:00:28.79" resultid="19724" heatid="19937" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="3555" points="437" reactiontime="+69" swimtime="00:01:13.83" resultid="19725" heatid="19974" lane="6" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="285006" swrid="4690799" athleteid="19744">
              <RESULTS>
                <RESULT eventid="3551" points="376" swimtime="00:00:33.29" resultid="19745" heatid="19850" lane="2" entrytime="00:00:32.50" />
                <RESULT eventid="3649" points="385" swimtime="00:02:20.17" resultid="19746" heatid="19894" lane="5" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="347" swimtime="00:00:29.75" resultid="19747" heatid="19953" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="3512" points="348" swimtime="00:02:39.05" resultid="19748" heatid="19999" lane="6" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="226836" swrid="4406865" athleteid="19749">
              <RESULTS>
                <RESULT eventid="9711" points="444" reactiontime="+90" swimtime="00:02:29.38" resultid="19750" heatid="19830" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="498" swimtime="00:00:26.37" resultid="19751" heatid="19958" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="3562" points="442" reactiontime="+75" swimtime="00:01:05.40" resultid="19752" heatid="19981" lane="6" entrytime="00:01:02.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="295252" swrid="4690789" athleteid="19769">
              <RESULTS>
                <RESULT eventid="3547" points="464" swimtime="00:00:34.93" resultid="19770" heatid="19843" lane="7" entrytime="00:00:34.50" />
                <RESULT eventid="3570" points="476" reactiontime="+73" swimtime="00:02:24.66" resultid="19771" heatid="19885" lane="2" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="465" swimtime="00:00:30.62" resultid="19772" heatid="19931" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="3505" points="433" swimtime="00:02:44.94" resultid="19773" heatid="19990" lane="6" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="285010" swrid="4690802" athleteid="19753">
              <RESULTS>
                <RESULT eventid="3628" points="351" reactiontime="+89" swimtime="00:01:23.04" resultid="19754" heatid="19871" lane="8" entrytime="00:01:19.00" />
                <RESULT eventid="3594" points="411" swimtime="00:00:28.12" resultid="19755" heatid="19953" lane="7" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="287369" swrid="4690795" athleteid="19736">
              <RESULTS>
                <RESULT eventid="3547" points="481" swimtime="00:00:34.53" resultid="19737" heatid="19843" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="3590" points="477" swimtime="00:00:30.36" resultid="19738" heatid="19932" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="3505" points="498" swimtime="00:02:37.42" resultid="19739" heatid="19991" lane="4" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="GER" license="266174" swrid="4558991" athleteid="19756">
              <RESULTS>
                <RESULT eventid="3547" points="569" swimtime="00:00:32.64" resultid="19757" heatid="19844" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="3570" points="572" reactiontime="+75" swimtime="00:02:16.08" resultid="19758" heatid="19888" lane="8" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="530" swimtime="00:00:29.31" resultid="19759" heatid="19935" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="3505" points="467" swimtime="00:02:40.81" resultid="19760" heatid="19992" lane="5" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="156716" swrid="4078097" athleteid="19761">
              <RESULTS>
                <RESULT eventid="3649" points="567" reactiontime="+65" swimtime="00:02:03.19" resultid="19762" heatid="19899" lane="3" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="532" swimtime="00:00:25.80" resultid="19763" heatid="19958" lane="3" entrytime="00:00:24.80" />
                <RESULT eventid="3562" points="492" reactiontime="+60" swimtime="00:01:03.07" resultid="19764" heatid="19982" lane="1" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="GER" license="226832" swrid="4320785" athleteid="19732">
              <RESULTS>
                <RESULT eventid="3628" points="398" reactiontime="+74" swimtime="00:01:19.63" resultid="19733" heatid="19871" lane="2" entrytime="00:01:16.00" />
                <RESULT eventid="3545" points="371" reactiontime="+82" swimtime="00:02:57.03" resultid="19734" heatid="19915" lane="7" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3594" points="379" swimtime="00:00:28.89" resultid="19735" heatid="19954" lane="2" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="12820" points="437" swimtime="00:04:33.04" resultid="19774" heatid="20141" lane="8" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="200" swimtime="00:02:32.68" />
                    <SPLIT distance="300" swimtime="00:03:37.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19744" number="1" />
                    <RELAYPOSITION athleteid="19732" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="19749" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="19761" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="3574" points="503" swimtime="00:04:51.95" resultid="19775" heatid="20139" lane="2" entrytime="00:04:47.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="200" swimtime="00:02:34.84" />
                    <SPLIT distance="300" swimtime="00:03:47.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19736" number="1" />
                    <RELAYPOSITION athleteid="19726" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="19721" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="19756" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="UNBR" nation="CZE" clubid="14059" swrid="73404" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="1994-01-01" firstname="Julia" gender="M" lastname="Janke-Frosch" nation="CZE" athleteid="17490">
              <RESULTS>
                <RESULT eventid="3551" points="616" swimtime="00:00:28.25" resultid="17491" heatid="19852" lane="2" entrytime="00:00:28.70" />
                <RESULT eventid="3649" points="568" reactiontime="+72" swimtime="00:02:03.15" resultid="17492" heatid="19899" lane="8" entrytime="00:02:00.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3562" points="621" reactiontime="+69" swimtime="00:00:58.38" resultid="17493" heatid="19982" lane="7" entrytime="00:00:59.70" />
                <RESULT eventid="3512" points="514" swimtime="00:02:19.66" resultid="17494" heatid="20001" lane="2" entrytime="00:02:18.60">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3605" points="582" swimtime="00:01:02.19" resultid="17495" heatid="20022" lane="6" entrytime="00:01:00.20" />
                <RESULT eventid="3613" points="594" swimtime="00:00:26.68" resultid="17496" heatid="20039" lane="1" entrytime="00:00:27.10" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STJO" nation="AUT" region="TLSV" clubid="14110" swrid="68105" name="Breedy Badger">
          <ATHLETES>
            <ATHLETE birthdate="2003-03-17" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43365" swrid="4826137" athleteid="18012">
              <RESULTS>
                <RESULT eventid="3639" points="297" reactiontime="+94" swimtime="00:03:08.99" resultid="18013" heatid="19811" lane="6" entrytime="00:03:15.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="234" reactiontime="+89" swimtime="00:01:44.54" resultid="18014" heatid="19855" lane="8" entrytime="00:01:43.79" entrycourse="LCM" />
                <RESULT eventid="3570" points="294" swimtime="00:02:49.76" resultid="18015" heatid="19880" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="293" swimtime="00:00:35.72" resultid="18016" heatid="19923" lane="2" entrytime="00:00:37.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-11" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="37374" swrid="4639773" athleteid="18027">
              <RESULTS>
                <RESULT eventid="3621" points="362" swimtime="00:01:30.35" resultid="18028" heatid="19859" lane="5" entrytime="00:01:29.63" entrycourse="LCM" />
                <RESULT eventid="3538" points="364" swimtime="00:03:16.12" resultid="18029" heatid="19906" lane="5" entrytime="00:03:27.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="376" swimtime="00:00:32.86" resultid="18030" heatid="19928" lane="5" entrytime="00:00:32.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-09-09" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="37373" swrid="4639772" athleteid="18022">
              <RESULTS>
                <RESULT eventid="3639" points="418" reactiontime="+68" swimtime="00:02:48.63" resultid="18023" heatid="19819" lane="2" entrytime="00:02:41.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="414" swimtime="00:01:26.45" resultid="18024" heatid="19860" lane="5" entrytime="00:01:26.22" entrycourse="LCM" />
                <RESULT eventid="3570" points="451" reactiontime="+66" swimtime="00:02:27.26" resultid="18025" heatid="19885" lane="4" entrytime="00:02:22.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="493" swimtime="00:00:30.03" resultid="18026" heatid="19933" lane="2" entrytime="00:00:30.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2005-09-13" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="43366" swrid="4826138" athleteid="18017">
              <RESULTS>
                <RESULT eventid="3621" points="190" swimtime="00:01:52.00" resultid="18018" heatid="19854" lane="3" entrytime="00:01:46.46" entrycourse="SCM" />
                <RESULT eventid="3570" points="182" reactiontime="+73" swimtime="00:03:19.03" resultid="18019" heatid="19876" lane="6" entrytime="00:03:05.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="257" swimtime="00:00:37.29" resultid="18020" heatid="19923" lane="6" entrytime="00:00:37.42" entrycourse="LCM" />
                <RESULT eventid="3547" points="211" swimtime="00:00:45.42" resultid="18021" heatid="19837" lane="3" entrytime="00:00:46.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-08-30" firstname="Julia" gender="F" lastname="Janke-Frosch" nation="AUT" license="41133" swrid="4826143" athleteid="18031">
              <RESULTS>
                <RESULT eventid="3639" points="378" reactiontime="+84" swimtime="00:02:54.32" resultid="18032" heatid="19816" lane="2" entrytime="00:02:54.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3621" points="385" reactiontime="+87" swimtime="00:01:28.58" resultid="18033" heatid="19860" lane="8" entrytime="00:01:28.95" entrycourse="LCM" />
                <RESULT eventid="3570" points="400" swimtime="00:02:33.32" resultid="18034" heatid="19882" lane="3" entrytime="00:02:31.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3590" points="470" swimtime="00:00:30.51" resultid="18035" heatid="19930" lane="1" entrytime="00:00:31.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="UNATTACHED">
          <ATHLETES>
            <ATHLETE gender="F" lastname="Janke-Frosch" athleteid="20201">
              <RESULTS>
                <RESULT eventid="15972" status="WDR" swimtime="00:00:00.00" resultid="20203" late="yes" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
